//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "Cubo-Piramide.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply1 w4;    //: /sn:0 {0}(218,33)(110,33){1}
//: {2}(108,31)(108,-18){3}
//: {4}(108,35)(108,53)(218,53){5}
supply0 w22;    //: /sn:0 {0}(1072,360)(1122,360)(1122,371){1}
reg [7:0] w0;    //: /sn:0 {0}(#:510,68)(510,54){1}
//: {2}(510,50)(#:510,12){3}
//: {4}(#:508,52)(422,52)(422,-51){5}
reg [7:0] w12;    //: /sn:0 {0}(#:706,83)(670,83)(670,46){1}
//: {2}(#:672,44)(747,44)(747,-52){3}
//: {4}(670,42)(#:670,7){5}
supply0 w1;    //: /sn:0 {0}(218,103)(55,103){1}
//: {2}(53,101)(53,95){3}
//: {4}(55,93)(218,93){5}
//: {6}(53,91)(53,63){7}
//: {8}(55,61)(62,61)(62,83)(218,83){9}
//: {10}(53,59)(53,45){11}
//: {12}(55,43)(69,43)(69,73)(218,73){13}
//: {14}(53,41)(53,19){15}
//: {16}(55,17)(77,17)(77,63)(218,63){17}
//: {18}(53,15)(53,-7){19}
//: {20}(55,-9)(85,-9)(85,43)(218,43){21}
//: {22}(53,-11)(53,-22)(28,-22)(28,-16){23}
//: {24}(53,105)(53,110){25}
reg w11;    //: /sn:0 {0}(299,720)(284,720)(284,688)(216,688){1}
reg w9;    //: /sn:0 {0}(468,94)(446,94)(446,133)(724,133){1}
//: {2}(728,133)(743,133)(743,112){3}
//: {4}(726,135)(726,509){5}
//: {6}(724,511)(676,511){7}
//: {8}(726,513)(726,731)(665,731){9}
//: {10}(661,731)(540,731){11}
//: {12}(536,731)(385,731)(385,635)(216,635){13}
//: {14}(538,733)(538,746){15}
//: {16}(663,733)(663,815){17}
//: {18}(665,817)(1344,817)(1344,549)(1321,549){19}
//: {20}(663,819)(663,880)(230,880)(230,834)(288,834){21}
wire [7:0] w13;    //: /sn:0 {0}(#:442,546)(442,621)(833,621)(833,505){1}
wire [7:0] w6;    //: /sn:0 {0}(#:414,355)(335,355)(335,356)(325,356){1}
//: {2}(#:321,356)(209,356)(209,342){3}
//: {4}(323,358)(323,375)(208,375)(208,392){5}
wire [3:0] w16;    //: /sn:0 {0}(#:83,577)(83,632){1}
//: {2}(85,634)(#:112,634){3}
//: {4}(81,634)(53,634)(53,530){5}
//: {6}(53,529)(53,445){7}
//: {8}(53,444)(53,394){9}
//: {10}(53,393)(53,292){11}
//: {12}(53,291)(#:53,259){13}
wire w7;    //: /sn:0 {0}(57,445)(120,445)(120,479)(277,479)(277,510)(414,510){1}
wire [7:0] w25;    //: /sn:0 {0}(#:1020,612)(1020,652)(1261,652){1}
//: {2}(1263,650)(#:1263,577){3}
//: {4}(1263,654)(1263,732)(1196,732)(1196,707){5}
wire [7:0] w3;    //: /sn:0 {0}(#:318,208)(318,131){1}
//: {2}(318,127)(318,98)(348,98)(348,19){3}
//: {4}(316,129)(256,129)(256,68)(#:224,68){5}
wire [7:0] w20;    //: /sn:0 {0}(#:1262,523)(1262,500){1}
//: {2}(#:1264,498)(1313,498)(1313,475){3}
//: {4}(1262,496)(1262,131)(1214,131)(#:1214,189){5}
wire w29;    //: /sn:0 {0}(945,576)(770,576)(770,700)(410,700)(410,600)(253,600)(253,530)(57,530){1}
wire [7:0] w18;    //: /sn:0 {0}(#:862,256)(862,299)(967,299)(#:967,330){1}
wire [7:0] w23;    //: /sn:0 {0}(#:999,545)(#:999,389){1}
wire [7:0] w10;    //: /sn:0 {0}(#:471,479)(#:471,385){1}
wire w24;    //: /sn:0 {0}(830,351)(830,359)(943,359){1}
wire w31;    //: /sn:0 {0}(57,292)(117,292)(117,240)(298,240){1}
wire [7:0] w32;    //: /sn:0 {0}(#:818,191)(818,135){1}
//: {2}(820,133)(1121,133)(#:1121,189){3}
//: {4}(818,131)(818,82)(#:783,82){5}
wire w8;    //: /sn:0 {0}(1101,221)(1038,221)(1038,97)(1413,97)(1413,916)(751,916){1}
//: {2}(749,914)(749,223)(798,223){3}
//: {4}(747,916)(-45,916)(-45,394)(48,394){5}
wire [7:0] w17;    //: /sn:0 {0}(#:508,323)(#:508,122){1}
wire [7:0] w27;    //: /sn:0 {0}(#:590,773)(615,773){1}
//: {2}(619,773)(971,773)(#:971,612){3}
//: {4}(617,775)(617,818){5}
wire [1:0] w28;    //: /sn:0 {0}(#:112,694)(30,694)(30,672){1}
wire [7:0] w14;    //: /sn:0 {0}(#:617,485)(617,451){1}
//: {2}(#:619,449)(670,449)(670,411){3}
//: {4}(617,447)(617,149)(911,149)(#:911,191){5}
wire [7:0] w2;    //: /sn:0 {0}(#:490,772)(436,772){1}
//: {2}(432,772)(-6,772)(-6,183)(411,183)(#:411,208){3}
//: {4}(434,774)(434,815){5}
wire [7:0] w15;    //: /sn:0 {0}(#:1165,254)(1165,292)(1043,292)(#:1043,330){1}
wire [7:0] w5;    //: /sn:0 {0}(#:362,273)(362,290)(438,290)(#:438,323){1}
wire [7:0] w26;    //: /sn:0 {0}(#:618,539)(618,576){1}
//: {2}(616,578)(494,578)(#:494,546){3}
//: {4}(618,580)(618,598)(668,598)(668,584){5}
//: enddecls

  //: frame g44 @(273,796) /sn:0 /wi:69 /ht:68 /tx:"CLOCK"
  //: joint g8 (w1) @(53, 17) /w:[ 16 18 -1 15 ]
  //: frame g4 @(13,-34) /sn:0 /wi:390 /ht:183 /tx:"COSTANTE = 5"
  //: joint g16 (w32) @(818, 133) /w:[ 2 4 -1 1 ]
  myDEMUX8x2 g47 (.in(w23), .c(w29), .out1(w27), .out2(w25));   //: @(946, 546) /sz:(106, 65) /R:3 /sn:0 /p:[ Ti0>0 Li0>0 Bo0<3 Bo1<0 ]
  //: joint g3 (w4) @(108, 33) /w:[ 1 2 -1 4 ]
  //: joint g26 (w3) @(318, 129) /w:[ -1 2 4 1 ]
  myMUL8 g17 (.A(w5), .B(w17), .Cout(w6), .out(w10));   //: @(416, 324) /sz:(118, 60) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<1 ]
  //: VDD g2 (w4) @(119,-18) /sn:0 /w:[ 3 ]
  myMUX8x2 g30 (.a(w32), .b(w14), .c(w8), .out(w18));   //: @(799, 192) /sz:(132, 63) /R:3 /sn:0 /p:[ Ti0>0 Ti1>5 Li0>3 Bo0<0 ]
  //: joint g23 (w16) @(83, 634) /w:[ 2 1 4 -1 ]
  //: joint g24 (w9) @(726, 133) /w:[ 2 -1 1 4 ]
  //: GROUND g39 (w22) @(1122,377) /sn:0 /w:[ 1 ]
  assign w3 = {w1, w1, w1, w1, w1, w4, w1, w4}; //: CONCAT g1  @(223,68) /sn:0 /w:[ 5 0 5 9 13 17 5 21 0 ] /dr:1 /tp:0 /drp:1
  myREG8 g29 (.in(w26), .Clk(w9), .out(w14));   //: @(565, 486) /sz:(110, 52) /R:1 /sn:0 /p:[ Bi0>0 Ri0>7 To0<0 ]
  //: LED g60 (w6) @(209,335) /sn:0 /w:[ 3 ] /type:0
  //: LED g51 (w2) @(434,822) /sn:0 /R:2 /w:[ 5 ] /type:3
  myMUX8x2 g18 (.a(w3), .b(w2), .c(w31), .out(w5));   //: @(299, 209) /sz:(132, 63) /R:3 /sn:0 /p:[ Ti0>0 Ti1>3 Li0>1 Bo0<0 ]
  //: LED g70 (w0) @(422,-58) /sn:0 /w:[ 5 ] /type:3
  //: frame g25 @(155,313) /sn:0 /wi:180 /ht:132 /tx:"OVERFLOW"
  //: LED g65 (w16) @(83,570) /sn:0 /w:[ 0 ] /type:1
  //: joint g10 (w1) @(53, 61) /w:[ 8 10 -1 7 ]
  //: SWITCH g64 (w11) @(317,720) /sn:0 /R:2 /w:[ 0 ] /st:1 /dn:1
  //: joint g49 (w25) @(1263, 652) /w:[ -1 2 1 4 ]
  //: joint g72 (w0) @(510, 52) /w:[ -1 2 4 1 ]
  //: joint g50 (w9) @(538, 731) /w:[ 11 -1 12 14 ]
  assign w29 = w16[0]; //: TAP g6 @(51,530) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  //: frame g68 @(267,659) /sn:0 /wi:87 /ht:90 /tx:"ENABLE"
  //: joint g35 (w1) @(53, 103) /w:[ 1 2 -1 24 ]
  //: joint g9 (w1) @(53, 43) /w:[ 12 14 -1 11 ]
  //: joint g7 (w1) @(53, -9) /w:[ 20 22 -1 19 ]
  //: joint g56 (w9) @(663, 731) /w:[ 9 -1 10 16 ]
  //: joint g58 (w12) @(670, 44) /w:[ 2 4 -1 1 ]
  //: joint g22 (w9) @(726, 511) /w:[ -1 5 6 8 ]
  myREG8 g59 (.Clk(w9), .in(w27), .out(w2));   //: @(492, 747) /sz:(98, 54) /R:2 /sn:0 /p:[ Ti0>15 Ri0>0 Lo0<0 ]
  //: frame g71 @(773,450) /sn:0 /wi:122 /ht:78 /tx:"** RISULTATO **"
  //: joint g31 (w14) @(617, 449) /w:[ 2 4 -1 1 ]
  assign w31 = w16[3]; //: TAP g67 @(51,292) /sn:0 /R:2 /w:[ 0 11 12 ] /ss:1
  myADD8 g36 (.A(w18), .B(w15), .Cin(w22), .Cout(w24), .S(w23));   //: @(944, 331) /sz:(127, 57) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  myMUX8x2 g33 (.a(w32), .b(w20), .c(w8), .out(w15));   //: @(1102, 190) /sz:(132, 63) /R:3 /sn:0 /p:[ Ti0>3 Ti1>5 Li0>0 Bo0<0 ]
  //: SWITCH g45 (w9) @(306,834) /sn:0 /R:2 /w:[ 21 ] /st:1 /dn:1
  //: LED g41 (w20) @(1313,468) /sn:0 /w:[ 3 ] /type:3
  //: LED g54 (w27) @(617,825) /sn:0 /R:2 /w:[ 5 ] /type:3
  //: frame g69 @(802,321) /sn:0 /wi:66 /ht:66 /tx:"OVERFLOW"
  myREG8 g52 (.in(w25), .Clk(w9), .out(w20));   //: @(1209, 524) /sz:(111, 52) /R:1 /sn:0 /p:[ Bi0>3 Ri0>19 To0<0 ]
  assign w8 = w16[2]; //: TAP g40 @(51,394) /sn:0 /R:2 /w:[ 5 9 10 ] /ss:0
  //: joint g42 (w8) @(749, 916) /w:[ 1 2 4 -1 ]
  //: LED g66 (w28) @(30,665) /sn:0 /w:[ 1 ] /type:2
  assign w7 = w16[1]; //: TAP g12 @(51,445) /sn:0 /R:2 /w:[ 0 7 8 ] /ss:1
  //: LED g28 (w14) @(670,404) /sn:0 /w:[ 3 ] /type:3
  //: LED g34 (w26) @(668,577) /sn:0 /w:[ 5 ] /type:3
  //: LED g46 (w25) @(1196,700) /sn:0 /w:[ 5 ] /type:3
  //: LED g57 (w12) @(747,-59) /sn:0 /w:[ 3 ] /type:3
  //: joint g11 (w1) @(53, 93) /w:[ 4 6 -1 3 ]
  //: DIP g14 (w0) @(510,2) /sn:0 /w:[ 3 ] /st:4 /dn:1
  //: GROUND g5 (w1) @(28,-10) /sn:0 /w:[ 23 ]
  myREG8 g19 (.in(w12), .Clk(w9), .out(w32));   //: @(707, 56) /sz:(75, 56) /sn:0 /p:[ Li0>0 Bi0>3 Ro0<5 ]
  //: frame g21 @(590,-37) /sn:0 /wi:143 /ht:65 /tx:"APOTEMA = A"
  //: joint g61 (w6) @(323, 356) /w:[ 1 -1 2 4 ]
  //: DIP g20 (w12) @(670,-3) /sn:0 /w:[ 5 ] /st:3 /dn:1
  myDEMUX8x2 g32 (.in(w10), .c(w7), .out1(w13), .out2(w26));   //: @(415, 480) /sz:(112, 65) /R:3 /sn:0 /p:[ Ti0>0 Li0>1 Bo0<0 Bo1<3 ]
  //: joint g63 (w9) @(663, 817) /w:[ 18 17 -1 20 ]
  //: frame g15 @(432,-34) /sn:0 /wi:144 /ht:68 /tx:"LATO CUBO = L"
  //: LED g0 (w3) @(348,12) /sn:0 /w:[ 3 ] /type:3
  //: joint g38 (w26) @(618, 578) /w:[ -1 1 2 4 ]
  //: joint g43 (w20) @(1262, 498) /w:[ 2 4 -1 1 ]
  //: LED g48 (w13) @(833,498) /sn:0 /w:[ 1 ] /type:3
  //: LED g27 (w6) @(208,399) /sn:0 /R:2 /w:[ 5 ] /type:3
  //: LED g37 (w24) @(830,344) /sn:0 /w:[ 0 ] /type:0
  ControlUnit g62 (.enable(w11), .clk(w9), .n_clk(w28), .control(w16));   //: @(113, 614) /sz:(102, 98) /sn:0 /p:[ Ri0>1 Ri1>13 Lo0<0 Lo1<3 ]
  //: joint g55 (w27) @(617, 773) /w:[ 2 -1 1 4 ]
  myREG8 g13 (.in(w0), .Clk(w9), .out(w17));   //: @(469, 69) /sz:(83, 52) /R:3 /sn:0 /p:[ Ti0>0 Li0>0 Bo0<1 ]
  //: joint g53 (w2) @(434, 772) /w:[ 1 -1 2 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin myXOR
module myXOR(out, B, A);
//: interface  /sz:(85, 111) /bd:[ Li0>A(20/111) Li1>B(84/111) Ro0<out(54/111) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(380,285)(354,285)(354,315)(153,315){1}
//: {2}(151,313)(151,219)(111,219){3}
//: {4}(151,317)(151,431)(199,431){5}
input A;    //: /sn:0 {0}(240,205)(203,205){1}
//: {2}(201,203)(201,137)(111,137){3}
//: {4}(201,207)(201,372)(383,372){5}
output out;    //: /sn:0 {0}(634,315)(696,315){1}
wire w6;    //: /sn:0 {0}(473,270)(506,270)(506,303)(550,303){1}
wire w3;    //: /sn:0 {0}(383,400)(354,400)(354,431)(282,431){1}
wire w1;    //: /sn:0 {0}(311,205)(337,205)(337,258)(380,258){1}
wire w8;    //: /sn:0 {0}(476,384)(506,384)(506,331)(550,331){1}
//: enddecls

  myNAND2 g4 (.a(w1), .b(B), .out(w6));   //: @(381, 243) /sz:(91, 54) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  myNAND2 g8 (.a(A), .b(w3), .out(w8));   //: @(384, 356) /sz:(91, 57) /sn:0 /p:[ Li0>5 Li1>0 Ro0<0 ]
  MyINV g3 (.in(A), .out(w1));   //: @(241, 182) /sz:(69, 47) /sn:0 /p:[ Li0>0 Ro0<0 ]
  //: OUT g2 (out) @(693,315) /sn:0 /w:[ 1 ]
  //: IN g1 (B) @(109,219) /sn:0 /w:[ 3 ]
  //: joint g6 (A) @(201, 205) /w:[ 1 2 -1 4 ]
  myNAND2 g7 (.a(w6), .b(w8), .out(out));   //: @(551, 287) /sz:(82, 57) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: joint g9 (B) @(151, 315) /w:[ 1 2 -1 4 ]
  MyINV g5 (.in(B), .out(w3));   //: @(200, 407) /sz:(81, 49) /sn:0 /p:[ Li0>5 Ro0<1 ]
  //: IN g0 (A) @(109,137) /sn:0 /w:[ 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin myFA
module myFA(S, Cin, B, A, Cout);
//: interface  /sz:(97, 88) /bd:[ Ti0>B(17/97) Ti1>A(77/97) Ri0>Cin(39/88) Lo0<Cout(41/88) Bo0<S(48/97) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input B;    //: /sn:0 {0}(435,582)(99,582)(99,155){1}
//: {2}(99,151)(99,144)(256,144){3}
//: {4}(97,153)(65,153){5}
input A;    //: /sn:0 {0}(435,551)(168,551)(168,114){1}
//: {2}(170,112)(256,112){3}
//: {4}(166,112)(65,112){5}
input Cin;    //: /sn:0 {0}(66,499)(257,499){1}
//: {2}(261,499)(354,499)(354,316)(444,316){3}
//: {4}(259,497)(259,175)(517,175){5}
output Cout;    //: /sn:0 {0}(805,432)(876,432){1}
output S;    //: /sn:0 {0}(612,161)(862,161){1}
wire w3;    //: /sn:0 {0}(444,286)(398,286)(398,148){1}
//: {2}(400,146)(517,146){3}
//: {4}(398,144)(398,129)(358,129){5}
wire w8;    //: /sn:0 {0}(694,449)(608,449)(608,564)(553,564){1}
wire w5;    //: /sn:0 {0}(556,299)(608,299)(608,420)(694,420){1}
//: enddecls

  //: OUT g4 (S) @(859,161) /sn:0 /w:[ 1 ]
  myNAND2 g8 (.a(w3), .b(Cin), .out(w5));   //: @(445, 269) /sz:(110, 60) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  //: IN g3 (Cin) @(64,499) /sn:0 /w:[ 0 ]
  //: IN g2 (B) @(63,153) /sn:0 /w:[ 5 ]
  //: IN g1 (A) @(63,112) /sn:0 /w:[ 5 ]
  myXOR g10 (.B(Cin), .A(w3), .out(S));   //: @(518, 137) /sz:(93, 51) /sn:0 /p:[ Li0>5 Li1>3 Ro0<0 ]
  myNAND2 g6 (.a(A), .b(B), .out(w8));   //: @(436, 532) /sz:(116, 64) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: joint g7 (A) @(168, 112) /w:[ 2 -1 4 1 ]
  myNAND2 g9 (.a(w5), .b(w8), .out(Cout));   //: @(695, 403) /sz:(109, 59) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  //: joint g12 (w3) @(398, 146) /w:[ 2 4 -1 1 ]
  //: OUT g5 (Cout) @(873,432) /sn:0 /w:[ 1 ]
  //: joint g11 (B) @(99, 153) /w:[ -1 2 4 1 ]
  myXOR g0 (.B(B), .A(A), .out(w3));   //: @(257, 102) /sz:(100, 56) /sn:0 /p:[ Li0>3 Li1>3 Ro0<5 ]
  //: joint g13 (Cin) @(259, 499) /w:[ 2 4 1 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin myFFDet
module myFFDet(Y, Clk, D, Y_n);
//: interface  /sz:(108, 80) /bd:[ Li0>D(18/80) Bi0>Clk(48/108) Ro0<Y(19/80) Ro1<Y_n(35/80) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input Clk;    //: /sn:0 {0}(114,364)(152,364){1}
//: {2}(156,364)(423,364)(423,324){3}
//: {4}(154,362)(154,307)(185,307){5}
output Y_n;    //: /sn:0 {0}(468,302)(540,302)(540,329)(555,329){1}
input D;    //: /sn:0 {0}(106,201)(221,201)(221,183)(236,183){1}
output Y;    //: /sn:0 {0}(468,274)(482,274)(482,286)(574,286){1}
wire w4;    //: /sn:0 {0}(315,203)(300,203){1}
wire w1;    //: /sn:0 {0}(265,305)(294,305)(294,251)(264,251)(264,221){1}
wire w2;    //: /sn:0 {0}(300,179)(350,179)(350,278)(389,278){1}
//: enddecls

  //: frame g8 @(365,239) /sn:0 /wi:143 /ht:111 /tx:"SLAVE"
  //: OUT g4 (Y) @(571,286) /sn:0 /w:[ 1 ]
  //: IN g3 (Clk) @(112,364) /sn:0 /w:[ 0 ]
  //: IN g2 (D) @(104,201) /sn:0 /w:[ 0 ]
  //: joint g1 (Clk) @(154, 364) /w:[ 2 4 1 -1 ]
  //: OUT g6 (Y_n) @(552,329) /sn:0 /w:[ 1 ]
  //: frame g7 @(207,149) /sn:0 /wi:128 /ht:95 /tx:"MASTER"
  myFFD g9 (.D(D), .Clk(w1), .Y(w2), .Y_n(w4));   //: @(237, 167) /sz:(62, 53) /sn:0 /p:[ Li0>1 Bi0>1 Ro0<0 Ro1<1 ]
  MyINV g5 (.in(Clk), .out(w1));   //: @(186, 284) /sz:(78, 46) /sn:0 /p:[ Li0>5 Ro0<0 ]
  myFFD g0 (.D(w2), .Clk(Clk), .Y(Y), .Y_n(Y_n));   //: @(390, 259) /sz:(77, 64) /sn:0 /p:[ Li0>1 Bi0>3 Ro0<0 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myLATCHSR
module myLATCHSR(y_n, y, s, r);
//: interface  /sz:(163, 125) /bd:[ Li0>s(24/125) Li1>r(93/125) Ro0<y(22/125) Ro1<y_n(38/125) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input r;    //: /sn:0 {0}(190,265)(106,265){1}
output y_n;    //: /sn:0 {0}(190,236)(165,236)(165,196)(388,196){1}
//: {2}(392,196)(421,196)(421,170)(472,170){3}
//: {4}(390,194)(390,109)(297,109){5}
output y;    //: /sn:0 {0}(201,126)(163,126)(163,162)(364,162)(364,248){1}
//: {2}(366,250)(409,250)(409,273)(475,273){3}
//: {4}(362,250)(283,250){5}
input s;    //: /sn:0 {0}(104,97)(201,97){1}
//: enddecls

  //: OUT g4 (y_n) @(469,170) /sn:0 /w:[ 3 ]
  //: joint g3 (y) @(364, 250) /w:[ 2 1 4 -1 ]
  //: OUT g2 (y) @(472,273) /sn:0 /w:[ 3 ]
  myNOR2 g1 (.a(y_n), .b(r), .out(y));   //: @(191, 226) /sz:(91, 52) /sn:0 /p:[ Li0>0 Li1>0 Ro0<5 ]
  //: IN g6 (s) @(102,97) /sn:0 /w:[ 0 ]
  //: IN g7 (r) @(104,265) /sn:0 /w:[ 1 ]
  //: joint g5 (y_n) @(390, 196) /w:[ 2 4 1 -1 ]
  myNOR2 g0 (.a(s), .b(y), .out(y_n));   //: @(202, 88) /sz:(94, 51) /sn:0 /p:[ Li0>1 Li1>0 Ro0<5 ]

endmodule
//: /netlistEnd

//: /netlistBegin myMUX2
module myMUX2(c, out, in1, in0);
//: interface  /sz:(154, 104) /bd:[ Li0>in1(76/104) Li1>in0(23/104) Bi0>c(77/154) Ro0<out(51/104) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in1;    //: /sn:0 {0}(142,341)(342,341)(342,439)(374,439){1}
input in0;    //: /sn:0 {0}(146,163)(338,163)(338,262)(364,262){1}
output out;    //: /sn:0 {0}(674,359)(735,359){1}
input c;    //: /sn:0 {0}(157,508)(196,508)(196,471){1}
//: {2}(198,469)(374,469){3}
//: {4}(196,467)(196,293)(221,293){5}
wire w7;    //: /sn:0 {0}(486,453)(522,453)(522,376)(564,376){1}
wire w4;    //: /sn:0 {0}(471,275)(521,275)(521,346)(564,346){1}
wire w1;    //: /sn:0 {0}(305,292)(364,292){1}
//: enddecls

  MyINV g4 (.in(c), .out(w1));   //: @(222, 266) /sz:(82, 53) /sn:0 /p:[ Li0>5 Ro0<0 ]
  //: joint g8 (c) @(196, 469) /w:[ 2 4 -1 1 ]
  //: IN g3 (c) @(155,508) /sn:0 /w:[ 0 ]
  //: OUT g2 (out) @(732,359) /sn:0 /w:[ 1 ]
  //: IN g1 (in1) @(140,341) /sn:0 /w:[ 0 ]
  myNAND2 g6 (.b(c), .a(in1), .out(w7));   //: @(375, 430) /sz:(110, 56) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  myNAND2 g7 (.b(w7), .a(w4), .out(out));   //: @(565, 337) /sz:(108, 55) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  myNAND2 g5 (.b(w1), .a(in0), .out(w4));   //: @(365, 252) /sz:(105, 57) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g0 (in0) @(144,163) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myREG8
module myREG8(Clk, out, in);
//: interface  /sz:(122, 206) /bd:[ Li0>in[7:0](102/206) Bi0>Clk(60/122) Ro0<out[7:0](99/206) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] in;    //: /sn:0 {0}(#:214,37)(332,37)(332,66){1}
//: {2}(332,67)(332,117){3}
//: {4}(332,118)(332,184)(332,184)(332,232){5}
//: {6}(332,233)(332,333){7}
//: {8}(332,334)(332,430){9}
//: {10}(332,431)(332,534){11}
//: {12}(332,535)(332,631){13}
//: {14}(332,632)(332,745){15}
//: {16}(332,746)(332,764){17}
input Clk;    //: /sn:0 {0}(454,475)(454,507)(307,507){1}
//: {2}(305,505)(305,450){3}
//: {4}(305,446)(305,389){5}
//: {6}(307,387)(454,387)(454,370){7}
//: {8}(305,385)(305,291){9}
//: {10}(307,289)(459,289)(459,265){11}
//: {12}(305,287)(305,195){13}
//: {14}(307,193)(458,193)(458,171){15}
//: {16}(305,191)(305,88)(457,88)(457,75){17}
//: {18}(303,448)(220,448){19}
//: {20}(305,509)(305,602){21}
//: {22}(307,604)(451,604)(451,579){23}
//: {24}(305,606)(305,711){25}
//: {26}(307,713)(446,713)(446,689){27}
//: {28}(305,715)(305,806)(444,806)(444,790){29}
output [7:0] out;    //: /sn:0 {0}(#:809,478)(938,478){1}
wire w6;    //: /sn:0 {0}(421,217)(371,217)(371,233)(336,233){1}
wire w13;    //: /sn:0 {0}(503,425)(597,425)(597,483)(803,483){1}
wire w16;    //: /sn:0 {0}(500,320)(615,320)(615,473)(803,473){1}
wire w7;    //: /sn:0 {0}(523,248)(508,248){1}
wire w4;    //: /sn:0 {0}(495,639)(554,639)(554,503)(803,503){1}
wire w0;    //: /sn:0 {0}(419,25)(373,25)(373,67)(336,67){1}
wire w3;    //: /sn:0 {0}(420,118)(336,118){1}
wire w22;    //: /sn:0 {0}(507,119)(687,119)(687,453)(803,453){1}
wire w20;    //: /sn:0 {0}(508,774)(493,774){1}
wire w12;    //: /sn:0 {0}(416,425)(362,425)(362,431)(336,431){1}
wire w18;    //: /sn:0 {0}(408,639)(383,639)(383,632)(336,632){1}
wire w19;    //: /sn:0 {0}(508,218)(656,218)(656,463)(803,463){1}
wire w23;    //: /sn:0 {0}(493,740)(583,740)(583,513)(803,513){1}
wire w10;    //: /sn:0 {0}(500,529)(521,529)(521,493)(803,493){1}
wire w21;    //: /sn:0 {0}(406,740)(366,740)(366,746)(336,746){1}
wire w1;    //: /sn:0 {0}(521,58)(506,58){1}
wire w8;    //: /sn:0 {0}(515,347)(500,347){1}
wire w17;    //: /sn:0 {0}(510,670)(495,670){1}
wire w14;    //: /sn:0 {0}(515,563)(500,563){1}
wire w2;    //: /sn:0 {0}(803,443)(736,443)(736,26)(506,26){1}
wire w11;    //: /sn:0 {0}(518,457)(503,457){1}
wire w15;    //: /sn:0 {0}(413,529)(379,529)(379,535)(336,535){1}
wire w5;    //: /sn:0 {0}(522,155)(507,155){1}
wire w9;    //: /sn:0 {0}(413,320)(354,320)(354,334)(336,334){1}
//: enddecls

  myFFDet g8 (.D(w12), .Clk(Clk), .Y_n(w11), .Y(w13));   //: @(417, 411) /sz:(85, 63) /sn:0 /p:[ Li0>0 Bi0>0 Ro0<1 Ro1<0 ]
  //: joint g4 (Clk) @(305, 193) /w:[ 14 16 -1 13 ]
  myFFDet g3 (.D(w0), .Clk(Clk), .Y_n(w1), .Y(w2));   //: @(420, 12) /sz:(85, 62) /sn:0 /p:[ Li0>0 Bi0>17 Ro0<1 Ro1<1 ]
  //: joint g16 (Clk) @(305, 604) /w:[ 22 21 -1 24 ]
  //: joint g17 (Clk) @(305, 507) /w:[ 1 2 -1 20 ]
  assign out = {w2, w22, w19, w16, w13, w10, w4, w23}; //: CONCAT g26  @(808,478) /sn:0 /w:[ 0 0 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  //: IN g2 (Clk) @(218,448) /sn:0 /w:[ 19 ]
  assign w15 = in[2]; //: TAP g23 @(330,535) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  //: OUT g1 (out) @(935,478) /sn:0 /w:[ 1 ]
  assign w18 = in[1]; //: TAP g24 @(330,632) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  assign w0 = in[7]; //: TAP g18 @(330,67) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  myFFDet g10 (.D(w18), .Clk(Clk), .Y_n(w17), .Y(w4));   //: @(409, 625) /sz:(85, 63) /sn:0 /p:[ Li0>0 Bi0>27 Ro0<1 Ro1<0 ]
  assign w21 = in[0]; //: TAP g25 @(330,746) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  myFFDet g6 (.D(w6), .Clk(Clk), .Y_n(w7), .Y(w19));   //: @(422, 204) /sz:(85, 60) /sn:0 /p:[ Li0>0 Bi0>11 Ro0<1 Ro1<0 ]
  myFFDet g7 (.D(w9), .Clk(Clk), .Y_n(w8), .Y(w16));   //: @(414, 306) /sz:(85, 63) /sn:0 /p:[ Li0>0 Bi0>7 Ro0<1 Ro1<0 ]
  myFFDet g9 (.D(w15), .Clk(Clk), .Y_n(w14), .Y(w10));   //: @(414, 515) /sz:(85, 63) /sn:0 /p:[ Li0>0 Bi0>23 Ro0<1 Ro1<0 ]
  assign w12 = in[3]; //: TAP g22 @(330,431) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  //: joint g12 (Clk) @(305, 289) /w:[ 10 12 -1 9 ]
  myFFDet g5 (.D(w3), .Clk(Clk), .Y_n(w5), .Y(w22));   //: @(421, 104) /sz:(85, 66) /sn:0 /p:[ Li0>0 Bi0>15 Ro0<1 Ro1<0 ]
  myFFDet g11 (.D(w21), .Clk(Clk), .Y_n(w20), .Y(w23));   //: @(407, 726) /sz:(85, 63) /sn:0 /p:[ Li0>0 Bi0>29 Ro0<1 Ro1<0 ]
  //: joint g14 (Clk) @(305, 448) /w:[ -1 4 18 3 ]
  assign w3 = in[6]; //: TAP g19 @(330,118) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  assign w9 = in[4]; //: TAP g21 @(330,334) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  assign w6 = in[5]; //: TAP g20 @(330,233) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  //: IN g0 (in) @(212,37) /sn:0 /w:[ 0 ]
  //: joint g15 (Clk) @(305, 713) /w:[ 26 25 -1 28 ]
  //: joint g13 (Clk) @(305, 387) /w:[ 6 8 -1 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin myAND2
module myAND2(out, b, a);
//: interface  /sz:(102, 81) /bd:[ Li0>a(13/81) Li1>b(63/81) Ro0<out(40/81) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(168,310)(231,310){1}
output out;    //: /sn:0 {0}(445,283)(487,283)(487,284)(493,284){1}
input a;    //: /sn:0 {0}(167,264)(231,264){1}
wire w0;    //: /sn:0 {0}(324,283)(352,283){1}
//: enddecls

  //: OUT g4 (out) @(490,284) /sn:0 /w:[ 1 ]
  //: IN g3 (b) @(166,310) /sn:0 /w:[ 0 ]
  //: IN g2 (a) @(165,264) /sn:0 /w:[ 0 ]
  MyINV g1 (.in(w0), .out(out));   //: @(353, 252) /sz:(91, 62) /sn:0 /p:[ Li0>1 Ro0<0 ]
  myNAND2 g0 (.b(b), .a(a), .out(w0));   //: @(232, 236) /sz:(91, 94) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myMUX8x2
module myMUX8x2(b, c, a, out);
//: interface  /sz:(126, 188) /bd:[ Li0>b[7:0](160/188) Li1>a[7:0](28/188) Bi0>c(63/126) Ro0<out[7:0](90/188) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] b;    //: /sn:0 {0}(#:236,775)(236,754){1}
//: {2}(236,753)(236,665){3}
//: {4}(236,664)(236,559){5}
//: {6}(236,558)(236,511)(237,511)(237,465){7}
//: {8}(237,464)(237,412)(236,412)(236,356){9}
//: {10}(236,355)(236,252){11}
//: {12}(236,251)(236,190){13}
//: {14}(236,189)(236,122){15}
//: {16}(236,121)(236,77)(#:65,77){17}
output [7:0] out;    //: /sn:0 {0}(#:743,345)(814,345){1}
input [7:0] a;    //: /sn:0 {0}(#:310,767)(310,732){1}
//: {2}(310,731)(310,631){3}
//: {4}(310,630)(310,531){5}
//: {6}(310,530)(310,437){7}
//: {8}(310,436)(310,386)(311,386)(311,325){9}
//: {10}(311,324)(311,222){11}
//: {12}(311,221)(311,142){13}
//: {14}(311,141)(311,68){15}
//: {16}(311,67)(311,30)(#:63,30){17}
input c;    //: /sn:0 {0}(526,674)(526,685)(134,685){1}
//: {2}(132,683)(132,599){3}
//: {4}(134,597)(527,597)(527,562){5}
//: {6}(132,595)(132,495){7}
//: {8}(134,493)(526,493)(526,461){9}
//: {10}(132,491)(132,394){11}
//: {12}(134,392)(522,392)(522,369){13}
//: {14}(132,390)(132,295){15}
//: {16}(134,293)(523,293)(523,271){17}
//: {18}(132,291)(132,205){19}
//: {20}(134,203)(523,203)(523,176){21}
//: {22}(132,201)(132,165){23}
//: {24}(134,163)(256,163)(256,133)(298,133)(298,104)(521,104)(521,73){25}
//: {26}(132,161)(132,140)(64,140){27}
//: {28}(132,687)(132,804)(528,804)(528,773){29}
wire w13;    //: /sn:0 {0}(466,326)(323,326)(323,325)(315,325){1}
wire w16;    //: /sn:0 {0}(470,445)(406,445)(406,465)(241,465){1}
wire w7;    //: /sn:0 {0}(737,320)(695,320)(695,147)(579,147){1}
wire w4;    //: /sn:0 {0}(467,160)(266,160)(266,190)(240,190){1}
wire w25;    //: /sn:0 {0}(470,631)(314,631){1}
wire w0;    //: /sn:0 {0}(465,30)(340,30)(340,68)(315,68){1}
wire w3;    //: /sn:0 {0}(577,44)(722,44)(722,310)(737,310){1}
wire w20;    //: /sn:0 {0}(471,546)(372,546)(372,559)(240,559){1}
wire w29;    //: /sn:0 {0}(471,730)(322,730)(322,732)(314,732){1}
wire w12;    //: /sn:0 {0}(466,353)(248,353)(248,356)(240,356){1}
wire w19;    //: /sn:0 {0}(737,350)(652,350)(652,432)(582,432){1}
wire w23;    //: /sn:0 {0}(737,360)(670,360)(670,533)(583,533){1}
wire w21;    //: /sn:0 {0}(471,519)(348,519)(348,531)(314,531){1}
wire w24;    //: /sn:0 {0}(470,658)(342,658)(342,665)(240,665){1}
wire w1;    //: /sn:0 {0}(465,57)(378,57)(378,87)(268,87)(268,122)(240,122){1}
wire w31;    //: /sn:0 {0}(737,380)(715,380)(715,744)(583,744){1}
wire w8;    //: /sn:0 {0}(467,255)(248,255)(248,252)(240,252){1}
wire w17;    //: /sn:0 {0}(470,418)(357,418)(357,437)(314,437){1}
wire w27;    //: /sn:0 {0}(737,370)(694,370)(694,645)(582,645){1}
wire w28;    //: /sn:0 {0}(471,757)(248,757)(248,754)(240,754){1}
wire w11;    //: /sn:0 {0}(737,330)(657,330)(657,242)(579,242){1}
wire w15;    //: /sn:0 {0}(737,340)(578,340){1}
wire w5;    //: /sn:0 {0}(467,133)(347,133)(347,142)(315,142){1}
wire w9;    //: /sn:0 {0}(467,228)(323,228)(323,222)(315,222){1}
//: enddecls

  myMUX2 g4 (.in1(w12), .in0(w13), .c(c), .out(w15));   //: @(467, 315) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>13 Ro0<1 ]
  myMUX2 g8 (.in1(w28), .in0(w29), .c(c), .out(w31));   //: @(472, 719) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>29 Ro0<1 ]
  myMUX2 g3 (.in1(w8), .in0(w9), .c(c), .out(w11));   //: @(468, 217) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>17 Ro0<1 ]
  assign w29 = a[7]; //: TAP g16 @(308,732) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  //: IN g17 (b) @(63,77) /sn:0 /w:[ 17 ]
  //: IN g26 (c) @(62,140) /sn:0 /w:[ 27 ]
  myMUX2 g2 (.in1(w4), .in0(w5), .c(c), .out(w7));   //: @(468, 122) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>21 Ro0<1 ]
  assign w20 = b[5]; //: TAP g23 @(234,559) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  //: joint g30 (c) @(132, 392) /w:[ 12 14 -1 11 ]
  //: IN g1 (a) @(61,30) /sn:0 /w:[ 17 ]
  assign w24 = b[6]; //: TAP g24 @(234,665) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  //: joint g29 (c) @(132, 293) /w:[ 16 18 -1 15 ]
  assign w1 = b[0]; //: TAP g18 @(234,122) /sn:0 /R:2 /w:[ 1 15 16 ] /ss:1
  assign w5 = a[1]; //: TAP g10 @(309,142) /sn:0 /R:2 /w:[ 1 13 14 ] /ss:1
  assign w28 = b[7]; //: TAP g25 @(234,754) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  myMUX2 g6 (.in1(w20), .in0(w21), .c(c), .out(w23));   //: @(472, 508) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>5 Ro0<1 ]
  myMUX2 g7 (.in1(w24), .in0(w25), .c(c), .out(w27));   //: @(471, 620) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>0 Ro0<1 ]
  assign w0 = a[0]; //: TAP g9 @(309,68) /sn:0 /R:2 /w:[ 1 15 16 ] /ss:1
  //: OUT g35 (out) @(811,345) /sn:0 /w:[ 1 ]
  assign w16 = b[4]; //: TAP g22 @(235,465) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  //: joint g31 (c) @(132, 493) /w:[ 8 10 -1 7 ]
  //: joint g33 (c) @(132, 685) /w:[ 1 2 -1 28 ]
  assign w13 = a[3]; //: TAP g12 @(309,325) /sn:0 /R:2 /w:[ 1 9 10 ] /ss:1
  //: joint g28 (c) @(132, 203) /w:[ 20 22 -1 19 ]
  assign out = {w31, w27, w23, w19, w15, w11, w7, w3}; //: CONCAT g34  @(742,345) /sn:0 /w:[ 0 0 0 0 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  myMUX2 g5 (.in1(w16), .in0(w17), .c(c), .out(w19));   //: @(471, 407) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>9 Ro0<1 ]
  assign w9 = a[2]; //: TAP g11 @(309,222) /sn:0 /R:2 /w:[ 1 11 12 ] /ss:1
  assign w21 = a[5]; //: TAP g14 @(308,531) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  assign w4 = b[1]; //: TAP g19 @(234,190) /sn:0 /R:2 /w:[ 1 13 14 ] /ss:1
  assign w12 = b[3]; //: TAP g21 @(234,356) /sn:0 /R:2 /w:[ 1 9 10 ] /ss:1
  assign w8 = b[2]; //: TAP g20 @(234,252) /sn:0 /R:2 /w:[ 1 11 12 ] /ss:1
  //: joint g32 (c) @(132, 597) /w:[ 4 6 -1 3 ]
  myMUX2 g0 (.in1(w1), .in0(w0), .c(c), .out(w3));   //: @(466, 19) /sz:(110, 53) /sn:0 /p:[ Li0>0 Li1>0 Bi0>25 Ro0<0 ]
  assign w25 = a[6]; //: TAP g15 @(308,631) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  //: joint g27 (c) @(132, 163) /w:[ 24 26 -1 23 ]
  assign w17 = a[4]; //: TAP g13 @(308,437) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin mySUMParziale
module mySUMParziale(B, A, out, s, Cout, Cin);
//: interface  /sz:(149, 113) /bd:[ Ti0>Cin(74/149) Li0>B[7:0](87/113) Li1>A[7:0](20/113) Bo0<Cout(74/149) Ro0<s(93/113) Ro1<out[7:0](54/113) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:41,103)(108,103){1}
//: {2}(109,103)(270,103){3}
//: {4}(271,103)(404,103){5}
//: {6}(405,103)(555,103){7}
//: {8}(556,103)(704,103){9}
//: {10}(705,103)(845,103){11}
//: {12}(846,103)(983,103){13}
//: {14}(984,103)(1139,103){15}
//: {16}(1140,103)(1183,103){17}
input [7:0] A;    //: /sn:0 {0}(#:41,65)(313,65){1}
//: {2}(314,65)(465,65){3}
//: {4}(466,65)(615,65){5}
//: {6}(616,65)(767,65){7}
//: {8}(768,65)(905,65){9}
//: {10}(906,65)(1042,65){11}
//: {12}(1043,65)(1216,65){13}
//: {14}(1217,65)(1297,65){15}
//: {16}(1298,65)(1332,65){17}
input Cin;    //: /sn:0 {0}(48,147)(169,147)(169,232){1}
output [7:0] out;    //: /sn:0 {0}(615,621)(#:615,521){1}
output Cout;    //: /sn:0 {0}(91,274)(59,274)(59,602)(324,602)(324,624){1}
output s;    //: /sn:0 {0}(1298,69)(1298,604)(1409,604){1}
wire w13;    //: /sn:0 {0}(630,515)(630,393)(878,393)(878,313){1}
wire w7;    //: /sn:0 {0}(970,263)(928,263){1}
wire w34;    //: /sn:0 {0}(109,232)(109,107){1}
wire w4;    //: /sn:0 {0}(1048,221)(1048,77)(1043,77)(1043,69){1}
wire w25;    //: /sn:0 {0}(462,229)(462,77)(466,77)(466,69){1}
wire w0;    //: /sn:0 {0}(1217,69)(1217,82)(1214,82)(1214,221){1}
wire w3;    //: /sn:0 {0}(1123,267)(1096,267)(1096,261)(1069,261){1}
wire w22;    //: /sn:0 {0}(535,269)(483,269){1}
wire w20;    //: /sn:0 {0}(613,227)(613,77)(616,77)(616,69){1}
wire w29;    //: /sn:0 {0}(260,231)(260,115)(271,115)(271,107){1}
wire w30;    //: /sn:0 {0}(320,231)(320,77)(314,77)(314,69){1}
wire w12;    //: /sn:0 {0}(829,265)(781,265){1}
wire w18;    //: /sn:0 {0}(620,515)(620,330)(731,330)(731,315){1}
wire w19;    //: /sn:0 {0}(553,227)(553,115)(556,115)(556,107){1}
wire w10;    //: /sn:0 {0}(907,223)(907,77)(906,77)(906,69){1}
wire w23;    //: /sn:0 {0}(610,515)(610,399)(585,399)(585,317){1}
wire w24;    //: /sn:0 {0}(402,229)(402,115)(405,115)(405,107){1}
wire w1;    //: /sn:0 {0}(1140,107)(1140,120)(1144,120)(1144,221){1}
wire w32;    //: /sn:0 {0}(242,273)(195,273)(195,272)(190,272){1}
wire w8;    //: /sn:0 {0}(1019,311)(1019,408)(640,408)(640,515){1}
wire w17;    //: /sn:0 {0}(682,267)(634,267){1}
wire w27;    //: /sn:0 {0}(384,271)(341,271){1}
wire w28;    //: /sn:0 {0}(600,515)(600,415)(433,415)(433,319){1}
wire w33;    //: /sn:0 {0}(590,515)(590,434)(291,434)(291,321){1}
wire w14;    //: /sn:0 {0}(700,225)(700,115)(705,115)(705,107){1}
wire w2;    //: /sn:0 {0}(1184,313)(1184,481)(650,481)(650,515){1}
wire w15;    //: /sn:0 {0}(760,225)(760,77)(768,77)(768,69){1}
wire w5;    //: /sn:0 {0}(988,221)(988,115)(984,115)(984,107){1}
wire w38;    //: /sn:0 {0}(580,515)(580,457)(140,457)(140,322){1}
wire w9;    //: /sn:0 {0}(847,223)(847,115)(846,115)(846,107){1}
//: enddecls

  myFA g4 (.B(w14), .A(w15), .Cin(w12), .Cout(w17), .S(w18));   //: @(683, 226) /sz:(97, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  myFA g8 (.B(w34), .A(Cin), .Cin(w32), .Cout(Cout), .S(w38));   //: @(92, 233) /sz:(97, 88) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: IN g16 (B) @(39,103) /sn:0 /w:[ 0 ]
  myFA g3 (.B(w9), .A(w10), .Cin(w7), .Cout(w12), .S(w13));   //: @(830, 224) /sz:(97, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w1 = B[0]; //: TAP g26 @(1140,101) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign s = A[0]; //: TAP g17 @(1298,63) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  //: IN g2 (A) @(39,65) /sn:0 /w:[ 0 ]
  //: OUT g30 (out) @(615,618) /sn:0 /R:3 /w:[ 0 ]
  assign w14 = B[3]; //: TAP g23 @(705,101) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign w9 = B[2]; //: TAP g24 @(846,101) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  myFA g1 (.B(w5), .A(w4), .Cin(w3), .Cout(w7), .S(w8));   //: @(971, 222) /sz:(97, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  assign out = {w38, w33, w28, w23, w18, w13, w8, w2}; //: CONCAT g29  @(615,520) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g18 (s) @(1406,604) /sn:0 /w:[ 1 ]
  assign w5 = B[1]; //: TAP g25 @(984,101) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  assign w25 = A[6]; //: TAP g10 @(466,63) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  myFA g6 (.B(w24), .A(w25), .Cin(w22), .Cout(w27), .S(w28));   //: @(385, 230) /sz:(97, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  myFA g7 (.B(w29), .A(w30), .Cin(w27), .Cout(w32), .S(w33));   //: @(243, 232) /sz:(97, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w30 = A[7]; //: TAP g9 @(314,63) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w19 = B[4]; //: TAP g22 @(556,101) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w15 = A[4]; //: TAP g12 @(768,63) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: OUT g28 (Cout) @(324,621) /sn:0 /R:3 /w:[ 1 ]
  myFA g5 (.B(w19), .A(w20), .Cin(w17), .Cout(w22), .S(w23));   //: @(536, 228) /sz:(97, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w20 = A[5]; //: TAP g11 @(616,63) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign w4 = A[2]; //: TAP g14 @(1043,63) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  assign w24 = B[5]; //: TAP g21 @(405,101) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign w34 = B[7]; //: TAP g19 @(109,101) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w29 = B[6]; //: TAP g20 @(271,101) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  myHA g0 (.b(w1), .a(w0), .out(w2), .cout(w3));   //: @(1124, 222) /sz:(110, 90) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bi0>0 Lo0<0 ]
  assign w0 = A[1]; //: TAP g15 @(1217,63) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  //: IN g27 (Cin) @(46,147) /sn:0 /w:[ 0 ]
  assign w10 = A[3]; //: TAP g13 @(906,63) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin myDEMUX8x2
module myDEMUX8x2(c, out2, in, out1);
//: interface  /sz:(144, 112) /bd:[ Li0>in[7:0](56/112) Bi0>c(68/144) Ro0<out1[7:0](27/112) Ro1<out2[7:0](79/112) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output [7:0] out2;    //: /sn:0 {0}(#:913,540)(1009,540){1}
input [7:0] in;    //: /sn:0 {0}(#:51,26)(163,26)(163,49){1}
//: {2}(163,50)(163,94)(164,94)(164,139){3}
//: {4}(164,140)(164,190)(163,190)(163,240){5}
//: {6}(163,241)(163,350){7}
//: {8}(163,351)(163,451){9}
//: {10}(163,452)(163,545){11}
//: {12}(163,546)(163,658){13}
//: {14}(163,659)(163,759){15}
//: {16}(163,760)(163,772){17}
output [7:0] out1;    //: /sn:0 {0}(#:909,412)(1000,412){1}
input c;    //: /sn:0 {0}(297,693)(297,711)(110,711){1}
//: {2}(108,709)(108,605){3}
//: {4}(110,603)(298,603)(298,588){5}
//: {6}(108,601)(108,511){7}
//: {8}(110,509)(301,509)(301,484){9}
//: {10}(108,507)(108,399){11}
//: {12}(110,397)(301,397)(301,378){13}
//: {14}(108,395)(108,302){15}
//: {16}(110,300)(299,300)(299,276){17}
//: {18}(108,298)(108,202){19}
//: {20}(110,200)(302,200)(302,180){21}
//: {22}(108,198)(108,103){23}
//: {24}(110,101)(301,101)(301,85){25}
//: {26}(108,99)(108,63)(48,63){27}
//: {28}(108,713)(108,807)(293,807)(293,796){29}
wire w16;    //: /sn:0 {0}(243,149)(176,149)(176,140)(168,140){1}
wire w34;    //: /sn:0 {0}(907,565)(590,565)(590,678)(363,678){1}
wire w39;    //: /sn:0 {0}(365,227)(434,227)(434,397)(903,397){1}
wire w36;    //: /sn:0 {0}(240,245)(175,245)(175,241)(167,241){1}
wire w22;    //: /sn:0 {0}(367,363)(693,363)(693,535)(907,535){1}
wire w20;    //: /sn:0 {0}(242,347)(191,347)(191,351)(167,351){1}
wire w30;    //: /sn:0 {0}(363,573)(540,573)(540,555)(907,555){1}
wire w42;    //: /sn:0 {0}(359,781)(640,781)(640,575)(907,575){1}
wire w19;    //: /sn:0 {0}(368,131)(456,131)(456,387)(903,387){1}
wire w18;    //: /sn:0 {0}(368,165)(766,165)(766,515)(907,515){1}
wire w12;    //: /sn:0 {0}(242,54)(175,54)(175,50)(167,50){1}
wire w23;    //: /sn:0 {0}(367,329)(473,329)(473,407)(903,407){1}
wire w24;    //: /sn:0 {0}(242,453)(222,453)(222,452)(167,452){1}
wire w31;    //: /sn:0 {0}(363,539)(510,539)(510,427)(903,427){1}
wire w32;    //: /sn:0 {0}(238,662)(175,662)(175,659)(167,659){1}
wire w27;    //: /sn:0 {0}(367,435)(490,435)(490,417)(903,417){1}
wire w35;    //: /sn:0 {0}(363,644)(533,644)(533,437)(903,437){1}
wire w28;    //: /sn:0 {0}(238,557)(175,557)(175,546)(167,546){1}
wire w14;    //: /sn:0 {0}(367,70)(796,70)(796,505)(907,505){1}
wire w15;    //: /sn:0 {0}(367,36)(574,36)(574,377)(903,377){1}
wire w38;    //: /sn:0 {0}(365,261)(745,261)(745,525)(907,525){1}
wire w43;    //: /sn:0 {0}(359,747)(583,747)(583,447)(903,447){1}
wire w26;    //: /sn:0 {0}(367,469)(666,469)(666,545)(907,545){1}
wire w40;    //: /sn:0 {0}(234,765)(175,765)(175,760)(167,760){1}
//: enddecls

  myDEMUX1x2 g8 (.in(w28), .c(c), .out2(w30), .out1(w31));   //: @(239, 530) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>5 Ro0<0 Ro1<0 ]
  myDEMUX1x2 g4 (.in(w12), .c(c), .out2(w14), .out1(w15));   //: @(243, 27) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>25 Ro0<0 Ro1<0 ]
  assign w36 = in[2]; //: TAP g3 @(161,241) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  assign w40 = in[7]; //: TAP g16 @(161,760) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  assign out2 = {w42, w34, w30, w26, w22, w38, w18, w14}; //: CONCAT g26  @(912,540) /sn:0 /w:[ 0 1 0 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: IN g17 (c) @(46,63) /sn:0 /w:[ 27 ]
  assign w16 = in[1]; //: TAP g2 @(162,140) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  //: joint g23 (c) @(108, 603) /w:[ 4 6 -1 3 ]
  //: joint g24 (c) @(108, 711) /w:[ 1 2 -1 28 ]
  assign w12 = in[0]; //: TAP g1 @(161,50) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: joint g18 (c) @(108, 101) /w:[ 24 26 -1 23 ]
  assign out1 = {w43, w35, w31, w27, w23, w39, w19, w15}; //: CONCAT g25  @(908,412) /sn:0 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  myDEMUX1x2 g10 (.in(w36), .c(c), .out2(w38), .out1(w39));   //: @(241, 218) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>17 Ro0<0 Ro1<0 ]
  myDEMUX1x2 g6 (.in(w20), .c(c), .out2(w22), .out1(w23));   //: @(243, 320) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>13 Ro0<0 Ro1<0 ]
  myDEMUX1x2 g9 (.in(w32), .c(c), .out2(w34), .out1(w35));   //: @(239, 635) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>0 Ro0<1 Ro1<0 ]
  myDEMUX1x2 g7 (.in(w24), .c(c), .out2(w26), .out1(w27));   //: @(243, 426) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>9 Ro0<0 Ro1<0 ]
  //: joint g22 (c) @(108, 509) /w:[ 8 10 -1 7 ]
  assign w20 = in[3]; //: TAP g12 @(161,351) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: OUT g28 (out2) @(1006,540) /sn:0 /w:[ 1 ]
  myDEMUX1x2 g11 (.in(w40), .c(c), .out2(w42), .out1(w43));   //: @(235, 738) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>29 Ro0<0 Ro1<0 ]
  myDEMUX1x2 g5 (.in(w16), .c(c), .out2(w18), .out1(w19));   //: @(244, 122) /sz:(123, 57) /sn:0 /p:[ Li0>0 Bi0>21 Ro0<0 Ro1<0 ]
  assign w28 = in[5]; //: TAP g14 @(161,546) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  //: joint g21 (c) @(108, 397) /w:[ 12 14 -1 11 ]
  //: joint g19 (c) @(108, 200) /w:[ 20 22 -1 19 ]
  //: joint g20 (c) @(108, 300) /w:[ 16 18 -1 15 ]
  //: IN g0 (in) @(49,26) /sn:0 /w:[ 0 ]
  assign w32 = in[6]; //: TAP g15 @(161,659) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  //: OUT g27 (out1) @(997,412) /sn:0 /w:[ 1 ]
  assign w24 = in[4]; //: TAP g13 @(161,452) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin myFFD
module myFFD(Y_n, D, Clk, Y);
//: interface  /sz:(107, 84) /bd:[ Li0>D(26/84) Bi0>Clk(47/107) Ro0<Y(20/84) Ro1<Y_n(36/84) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input Clk;    //: /sn:0 {0}(109,268)(389,268)(389,179){1}
output Y_n;    //: /sn:0 {0}(445,164)(478,164)(478,214)(532,214){1}
input D;    //: /sn:0 {0}(344,124)(143,124)(143,195){1}
//: {2}(145,197)(200,197){3}
//: {4}(141,197)(95,197){5}
output Y;    //: /sn:0 {0}(445,124)(492,124)(492,152)(560,152){1}
wire w0;    //: /sn:0 {0}(344,154)(312,154)(312,197)(287,197){1}
//: enddecls

  //: OUT g4 (Y_n) @(529,214) /sn:0 /w:[ 1 ]
  //: IN g3 (D) @(93,197) /sn:0 /w:[ 5 ]
  //: IN g2 (Clk) @(107,268) /sn:0 /w:[ 0 ]
  MyINV g1 (.in(D), .out(w0));   //: @(201, 174) /sz:(85, 47) /sn:0 /p:[ Li0>3 Ro0<1 ]
  myFFSR g7 (.S(D), .R(w0), .Clk(Clk), .Y(Y), .Y_n(Y_n));   //: @(345, 102) /sz:(99, 76) /sn:0 /p:[ Li0>0 Li1>0 Bi0>1 Ro0<0 Ro1<0 ]
  //: OUT g5 (Y) @(557,152) /sn:0 /w:[ 1 ]
  //: joint g0 (D) @(143, 197) /w:[ 2 1 4 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin myMUL8
module myMUL8(Cout, out, B, A);
//: interface  /sz:(86, 149) /bd:[ Li0>B[7:0](117/149) Li1>A[7:0](28/149) Bo0<Cout[7:0](45/86) Ro0<out[7:0](71/149) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:64,-18)(64,47){1}
//: {2}(64,48)(64,138){3}
//: {4}(64,139)(64,183)(63,183)(63,227){5}
//: {6}(63,228)(63,265)(64,265)(64,303){7}
//: {8}(64,304)(64,390){9}
//: {10}(64,391)(64,475){11}
//: {12}(64,476)(64,577){13}
//: {14}(64,578)(64,674){15}
//: {16}(64,675)(64,706){17}
input [7:0] A;    //: /sn:0 {0}(#:144,542)(44,542)(44,544)(34,544){1}
//: {2}(32,542)(32,446){3}
//: {4}(34,444)(44,444)(44,443)(#:141,443){5}
//: {6}(32,442)(32,359){7}
//: {8}(34,357)(44,357)(44,361)(#:141,361){9}
//: {10}(32,355)(32,277){11}
//: {12}(34,275)(#:140,275){13}
//: {14}(32,273)(32,187){15}
//: {16}(34,185)(44,185)(44,182)(#:139,182){17}
//: {18}(32,183)(32,107){19}
//: {20}(34,105)(112,105)(112,97)(#:140,97){21}
//: {22}(32,103)(32,15){23}
//: {24}(34,13)(46,13)(46,3)(101,3)(101,11)(#:142,11){25}
//: {26}(32,11)(#:32,-16){27}
//: {28}(32,546)(32,639)(#:145,639){29}
supply0 w0;    //: /sn:0 {0}(417,-12)(417,-33)(601,-33)(601,-5){1}
output [7:0] out;    //: /sn:0 {0}(801,-15)(801,33)(#:868,33)(#:868,52){1}
output [7:0] Cout;    //: /sn:0 {0}(#:1292,37)(1292,9)(865,9)(865,-12){1}
wire w6;    //: /sn:0 {0}(139,218)(75,218)(75,228)(67,228){1}
wire [7:0] w58;    //: /sn:0 {0}(#:1023,583)(1047,583)(1047,642)(930,642)(930,676)(#:941,676){1}
wire w50;    //: /sn:0 {0}(1297,43)(1297,231)(1216,231){1}
wire [7:0] w34;    //: /sn:0 {0}(#:596,129)(629,129)(629,179)(543,179)(543,216)(#:570,216){1}
wire w25;    //: /sn:0 {0}(892,492)(1009,492)(1009,240)(873,240)(873,58){1}
wire w39;    //: /sn:0 {0}(645,274)(645,311)(757,311)(757,324){1}
wire w3;    //: /sn:0 {0}(140,133)(76,133)(76,139)(68,139){1}
wire [7:0] w20;    //: /sn:0 {0}(#:285,560)(681,560)(681,604)(#:872,604){1}
wire [7:0] w29;    //: /sn:0 {0}(#:493,21)(520,21)(520,71)(435,71)(435,109)(#:445,109){1}
wire w42;    //: /sn:0 {0}(903,58)(903,195)(1013,195)(1013,68){1}
wire w18;    //: /sn:0 {0}(144,578)(68,578){1}
wire w12;    //: /sn:0 {0}(141,394)(76,394)(76,391)(68,391){1}
wire w63;    //: /sn:0 {0}(1327,43)(1327,757)(1016,757)(1016,734){1}
wire [7:0] w23;    //: /sn:0 {0}(#:286,657)(584,657)(584,717)(#:941,717){1}
wire w54;    //: /sn:0 {0}(1307,43)(1307,265)(1216,265){1}
wire w21;    //: /sn:0 {0}(145,675)(68,675){1}
wire w31;    //: /sn:0 {0}(1092,720)(1114,720)(1114,207)(893,207)(893,58){1}
wire w1;    //: /sn:0 {0}(142,45)(76,45)(76,48)(68,48){1}
wire [7:0] w32;    //: /sn:0 {0}(#:1092,696)(1212,696)(1212,292){1}
//: {2}(1212,291)(1212,265){3}
//: {4}(1212,264)(1212,231){5}
//: {6}(1212,230)(1212,216)(1211,216)(1211,203){7}
//: {8}(1211,202)(1211,181){9}
//: {10}(1211,180)(1211,162){11}
//: {12}(1211,161)(1211,119){13}
//: {14}(1211,118)(1211,64)(1013,64){15}
//: {16}(1012,64)(993,64){17}
wire [7:0] w46;    //: /sn:0 {0}(#:833,357)(849,357)(849,416)(705,416)(705,448)(#:741,448){1}
wire [7:0] w8;    //: /sn:0 {0}(#:280,200)(430,200)(430,150)(#:445,150){1}
wire [7:0] w52;    //: /sn:0 {0}(#:892,468)(918,468)(918,523)(845,523)(845,563)(#:872,563){1}
wire w44;    //: /sn:0 {0}(1215,162)(1267,162)(1267,43){1}
wire w27;    //: /sn:0 {0}(417,59)(417,81)(520,81)(520,96){1}
wire [7:0] w17;    //: /sn:0 {0}(#:282,461)(565,461)(565,489)(#:741,489){1}
wire w35;    //: /sn:0 {0}(596,153)(843,153)(843,58){1}
wire w33;    //: /sn:0 {0}(520,167)(520,191)(645,191)(645,203){1}
wire w28;    //: /sn:0 {0}(493,45)(769,45)(769,76)(833,76)(833,58){1}
wire w49;    //: /sn:0 {0}(1287,43)(1287,203)(1215,203){1}
wire w45;    //: /sn:0 {0}(757,395)(757,408)(816,408)(816,435){1}
wire [7:0] w14;    //: /sn:0 {0}(#:282,378)(#:682,378){1}
wire w48;    //: /sn:0 {0}(1277,43)(1277,181)(1215,181){1}
wire w41;    //: /sn:0 {0}(721,260)(853,260)(853,58){1}
wire [7:0] w11;    //: /sn:0 {0}(#:281,291)(555,291)(555,257)(#:570,257){1}
wire [7:0] w2;    //: /sn:0 {0}(#:283,28)(314,28)(314,1)(#:342,1){1}
wire w47;    //: /sn:0 {0}(863,58)(863,254)(961,254)(961,381)(833,381){1}
wire w15;    //: /sn:0 {0}(141,479)(76,479)(76,476)(68,476){1}
wire w55;    //: /sn:0 {0}(1317,43)(1317,292)(1216,292){1}
wire [7:0] w5;    //: /sn:0 {0}(#:281,115)(333,115)(333,42)(#:342,42){1}
wire w43;    //: /sn:0 {0}(1215,119)(1257,119)(1257,43){1}
wire w26;    //: /sn:0 {0}(1023,607)(1076,607)(1076,221)(883,221)(883,58){1}
wire w9;    //: /sn:0 {0}(140,307)(76,307)(76,304)(68,304){1}
wire w57;    //: /sn:0 {0}(947,621)(947,631)(1016,631)(1016,663){1}
wire w51;    //: /sn:0 {0}(816,506)(816,535)(947,535)(947,550){1}
wire [7:0] w40;    //: /sn:0 {0}(#:721,236)(737,236)(737,298)(661,298)(661,337)(#:682,337){1}
//: enddecls

  myPrParziale8 g8 (.m(w21), .M(A), .out(w23));   //: @(146, 627) /sz:(139, 62) /sn:0 /p:[ Li0>0 Li1>29 Ro0<0 ]
  myPrParziale8 g4 (.m(w9), .M(A), .out(w11));   //: @(141, 265) /sz:(139, 55) /sn:0 /p:[ Li0>0 Li1>13 Ro0<0 ]
  //: GROUND g44 (w0) @(601,1) /sn:0 /w:[ 1 ]
  assign Cout = {w63, w55, w54, w50, w49, w48, w44, w43}; //: CONCAT g16  @(1292,38) /sn:0 /R:1 /w:[ 0 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  myPrParziale8 g3 (.m(w6), .M(A), .out(w8));   //: @(140, 170) /sz:(139, 62) /sn:0 /p:[ Li0>0 Li1>17 Ro0<0 ]
  //: OUT g26 (Cout) @(865,-9) /sn:0 /R:1 /w:[ 1 ]
  assign w43 = w32[1]; //: TAP g17 @(1209,119) /sn:0 /R:2 /w:[ 0 13 14 ] /ss:1
  myPrParziale8 g2 (.m(w3), .M(A), .out(w5));   //: @(141, 85) /sz:(139, 62) /sn:0 /p:[ Li0>0 Li1>21 Ro0<0 ]
  assign w55 = w32[7]; //: TAP g23 @(1210,292) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:1
  //: joint g30 (A) @(32, 185) /w:[ 16 18 -1 15 ]
  assign w42 = w32[0]; //: TAP g24 @(1013,62) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  mySUMParziale g1 (.Cin(w0), .A(w2), .B(w5), .Cout(w27), .out(w29), .s(w28));   //: @(343, -11) /sz:(149, 69) /sn:0 /p:[ Ti0>0 Li0>1 Li1>1 Bo0<0 Ro0<0 Ro1<0 ]
  assign w9 = B[3]; //: TAP g39 @(62,304) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: joint g29 (A) @(32, 105) /w:[ 20 22 -1 19 ]
  assign w44 = w32[2]; //: TAP g18 @(1209,162) /sn:0 /R:2 /w:[ 0 11 12 ] /ss:1
  //: OUT g25 (out) @(801,-12) /sn:0 /R:1 /w:[ 0 ]
  mySUMParziale g10 (.Cin(w27), .A(w29), .B(w8), .Cout(w33), .out(w34), .s(w35));   //: @(446, 97) /sz:(149, 69) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<0 Ro0<0 Ro1<0 ]
  myPrParziale8 g6 (.m(w15), .M(A), .out(w17));   //: @(142, 431) /sz:(139, 62) /sn:0 /p:[ Li0>0 Li1>5 Ro0<0 ]
  assign out = {w42, w31, w26, w25, w47, w41, w35, w28}; //: CONCAT g9  @(868,53) /sn:0 /R:1 /w:[ 1 0 1 1 1 0 1 1 1 ] /dr:1 /tp:0 /drp:1
  myPrParziale8 g7 (.m(w18), .M(A), .out(w20));   //: @(145, 530) /sz:(139, 62) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: IN g35 (B) @(64,-20) /sn:0 /R:3 /w:[ 0 ]
  assign w48 = w32[3]; //: TAP g22 @(1209,181) /sn:0 /R:2 /w:[ 1 9 10 ] /ss:1
  //: joint g31 (A) @(32, 275) /w:[ 12 14 -1 11 ]
  //: joint g33 (A) @(32, 444) /w:[ 4 6 -1 3 ]
  assign w1 = B[0]; //: TAP g36 @(62,48) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  assign w15 = B[5]; //: TAP g41 @(62,476) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  assign w12 = B[4]; //: TAP g40 @(62,391) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  assign w21 = B[7]; //: TAP g42 @(62,675) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  mySUMParziale g12 (.Cin(w39), .A(w40), .B(w14), .Cout(w45), .out(w46), .s(w47));   //: @(683, 325) /sz:(149, 69) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<0 Ro0<0 Ro1<1 ]
  //: joint g28 (A) @(32, 13) /w:[ 24 26 -1 23 ]
  //: joint g34 (A) @(32, 544) /w:[ 1 2 -1 28 ]
  mySUMParziale g14 (.Cin(w51), .A(w52), .B(w20), .Cout(w57), .out(w58), .s(w26));   //: @(873, 551) /sz:(149, 69) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<0 Ro0<0 Ro1<0 ]
  mySUMParziale g11 (.Cin(w33), .A(w34), .B(w11), .Cout(w39), .out(w40), .s(w41));   //: @(571, 204) /sz:(149, 69) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<0 Ro0<0 Ro1<0 ]
  myPrParziale8 g5 (.m(w12), .M(A), .out(w14));   //: @(142, 350) /sz:(139, 58) /sn:0 /p:[ Li0>0 Li1>9 Ro0<0 ]
  assign w54 = w32[6]; //: TAP g21 @(1210,265) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  assign w49 = w32[4]; //: TAP g19 @(1209,203) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1
  assign w50 = w32[5]; //: TAP g20 @(1210,231) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  //: joint g32 (A) @(32, 357) /w:[ 8 10 -1 7 ]
  mySUMParziale g15 (.Cin(w57), .A(w58), .B(w23), .Cout(w63), .out(w32), .s(w31));   //: @(942, 664) /sz:(149, 69) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<1 Ro0<0 Ro1<0 ]
  myPrParziale8 g0 (.m(w1), .M(A), .out(w2));   //: @(143, 0) /sz:(139, 59) /sn:0 /p:[ Li0>0 Li1>25 Ro0<0 ]
  assign w6 = B[2]; //: TAP g38 @(61,228) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  assign w18 = B[6]; //: TAP g43 @(62,578) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  //: IN g27 (A) @(32,-18) /sn:0 /R:3 /w:[ 27 ]
  assign w3 = B[1]; //: TAP g37 @(62,139) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  mySUMParziale g13 (.Cin(w45), .A(w46), .B(w17), .Cout(w51), .out(w52), .s(w25));   //: @(742, 436) /sz:(149, 69) /sn:0 /p:[ Ti0>1 Li0>1 Li1>1 Bo0<0 Ro0<0 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myDEMUX1x2
module myDEMUX1x2(out2, out1, c, in);
//: interface  /sz:(123, 146) /bd:[ Li0>in(70/146) Bi0>c(58/123) Ro0<out2(112/146) Ro1<out1(25/146) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output out2;    //: /sn:0 {0}(432,440)(490,440)(490,378)(567,378){1}
input in;    //: /sn:0 {0}(337,423)(294,423)(294,235){1}
//: {2}(296,233)(319,233)(319,258)(341,258){3}
//: {4}(292,233)(73,233){5}
output out1;    //: /sn:0 {0}(431,274)(490,274)(490,329)(575,329){1}
input c;    //: /sn:0 {0}(337,455)(124,455)(124,409){1}
//: {2}(124,405)(124,288)(158,288){3}
//: {4}(122,407)(69,407){5}
wire w1;    //: /sn:0 {0}(249,288)(341,288){1}
//: enddecls

  //: joint g8 (c) @(124, 407) /w:[ -1 2 4 1 ]
  //: OUT g4 (out2) @(564,378) /sn:0 /w:[ 1 ]
  //: OUT g3 (out1) @(572,329) /sn:0 /w:[ 1 ]
  myAND2 g2 (.b(c), .a(in), .out(out2));   //: @(338, 415) /sz:(93, 52) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  myAND2 g1 (.b(w1), .a(in), .out(out1));   //: @(342, 250) /sz:(88, 50) /sn:0 /p:[ Li0>1 Li1>3 Ro0<0 ]
  //: IN g6 (c) @(67,407) /sn:0 /w:[ 5 ]
  //: joint g7 (in) @(294, 233) /w:[ 2 -1 4 1 ]
  //: IN g5 (in) @(71,233) /sn:0 /w:[ 5 ]
  MyINV g0 (.in(c), .out(w1));   //: @(159, 267) /sz:(89, 43) /sn:0 /p:[ Li0>3 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNOR2
module myNOR2(out, b, a);
//: interface  /sz:(141, 109) /bd:[ Li0>a(21/109) Li1>b(82/109) Ro0<out(46/109) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(288,265)(320,265){1}
//: {2}(324,265)(418,265)(418,290)(512,290){3}
//: {4}(322,267)(322,447)(553,447){5}
supply1 w0;    //: /sn:0 {0}(526,138)(526,202){1}
supply0 w1;    //: /sn:0 {0}(525,535)(525,487){1}
//: {2}(527,485)(567,485)(567,456){3}
//: {4}(523,485)(487,485)(487,419){5}
output out;    //: /sn:0 {0}(526,299)(526,332){1}
//: {2}(528,334)(643,334){3}
//: {4}(526,336)(526,384){5}
//: {6}(528,386)(567,386)(567,439){7}
//: {8}(524,386)(487,386)(487,402){9}
input a;    //: /sn:0 {0}(287,210)(378,210){1}
//: {2}(382,210)(512,210){3}
//: {4}(380,212)(380,410)(473,410){5}
wire w2;    //: /sn:0 {0}(526,219)(526,282){1}
//: enddecls

  _GGNMOS #(2, 1) g8 (.Z(out), .S(w1), .G(b));   //: @(561,447) /sn:0 /w:[ 7 3 5 ]
  //: GROUND g4 (w1) @(525,541) /sn:0 /w:[ 0 ]
  //: VDD g3 (w0) @(537,138) /sn:0 /w:[ 0 ]
  //: OUT g2 (out) @(640,334) /sn:0 /w:[ 3 ]
  //: IN g1 (b) @(286,265) /sn:0 /w:[ 0 ]
  //: joint g10 (out) @(526, 386) /w:[ 6 5 8 -1 ]
  _GGPMOS #(2, 1) g6 (.Z(out), .S(w2), .G(b));   //: @(520,290) /sn:0 /w:[ 0 1 3 ]
  //: joint g9 (w1) @(525, 485) /w:[ 2 -1 4 1 ]
  _GGNMOS #(2, 1) g7 (.Z(out), .S(w1), .G(a));   //: @(481,410) /sn:0 /w:[ 9 5 5 ]
  //: joint g12 (a) @(380, 210) /w:[ 2 -1 1 4 ]
  //: joint g11 (b) @(322, 265) /w:[ 2 -1 1 4 ]
  _GGPMOS #(2, 1) g5 (.Z(w2), .S(w0), .G(a));   //: @(520,210) /sn:0 /w:[ 0 1 3 ]
  //: IN g0 (a) @(285,210) /sn:0 /w:[ 0 ]
  //: joint g13 (out) @(526, 334) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNAND2
module myNAND2(out, b, a);
//: interface  /sz:(116, 124) /bd:[ Li0>a(37/124) Li1>b(98/124) Ro0<out(62/124) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(134,312)(229,312){1}
//: {2}(231,310)(231,195)(385,195){3}
//: {4}(231,314)(231,393)(349,393){5}
supply1 w0;    //: /sn:0 {0}(357,68)(357,131){1}
//: {2}(359,133)(399,133)(399,187){3}
//: {4}(355,133)(317,133)(317,145){5}
supply0 w1;    //: /sn:0 {0}(363,462)(363,402){1}
output out;    //: /sn:0 {0}(363,296)(363,266){1}
//: {2}(365,264)(479,264){3}
//: {4}(363,262)(363,218){5}
//: {6}(365,216)(399,216)(399,204){7}
//: {8}(361,216)(317,216)(317,162){9}
input a;    //: /sn:0 {0}(126,175)(280,175){1}
//: {2}(282,173)(282,153)(303,153){3}
//: {4}(282,177)(282,304)(349,304){5}
wire w2;    //: /sn:0 {0}(363,385)(363,313){1}
//: enddecls

  _GGNMOS #(2, 1) g8 (.Z(w2), .S(w1), .G(b));   //: @(357,393) /sn:0 /w:[ 0 1 5 ]
  //: GROUND g4 (w1) @(363,468) /sn:0 /w:[ 0 ]
  //: VDD g3 (w0) @(368,68) /sn:0 /w:[ 0 ]
  //: OUT g2 (out) @(476,264) /sn:0 /w:[ 3 ]
  //: IN g1 (b) @(132,312) /sn:0 /w:[ 0 ]
  //: joint g10 (out) @(363, 216) /w:[ 6 -1 8 5 ]
  _GGPMOS #(2, 1) g6 (.Z(out), .S(w0), .G(b));   //: @(393,195) /sn:0 /w:[ 7 3 3 ]
  //: joint g9 (w0) @(357, 133) /w:[ 2 1 4 -1 ]
  _GGNMOS #(2, 1) g7 (.Z(out), .S(w2), .G(a));   //: @(357,304) /sn:0 /w:[ 0 1 5 ]
  //: joint g12 (b) @(231, 312) /w:[ -1 2 1 4 ]
  //: joint g11 (a) @(282, 175) /w:[ -1 2 1 4 ]
  _GGPMOS #(2, 1) g5 (.Z(out), .S(w0), .G(a));   //: @(311,153) /sn:0 /w:[ 9 5 3 ]
  //: IN g0 (a) @(124,175) /sn:0 /w:[ 0 ]
  //: joint g13 (out) @(363, 264) /w:[ 2 4 -1 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin myFFSR
module myFFSR(Clk, R, Y, S, Y_n);
//: interface  /sz:(115, 93) /bd:[ Li0>S(27/93) Li1>R(64/93) Bi0>Clk(52/115) Ro0<Y(27/93) Ro1<Y_n(43/93) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input Clk;    //: /sn:0 {0}(95,266)(167,266){1}
//: {2}(169,264)(169,188)(210,188){3}
//: {4}(169,268)(169,328)(206,328){5}
input R;    //: /sn:0 {0}(85,359)(206,359){1}
output Y_n;    //: /sn:0 {0}(476,276)(499,276)(499,322)(556,322){1}
input S;    //: /sn:0 {0}(91,159)(210,159){1}
output Y;    //: /sn:0 {0}(583,275)(509,275)(509,244)(476,244){1}
wire w0;    //: /sn:0 {0}(297,345)(337,345)(337,277)(370,277){1}
wire w2;    //: /sn:0 {0}(297,175)(333,175)(333,245)(370,245){1}
//: enddecls

  //: joint g4 (Clk) @(169, 266) /w:[ -1 2 1 4 ]
  myLATCHSR g8 (.s(w2), .r(w0), .y(Y), .y_n(Y_n));   //: @(371, 234) /sz:(104, 59) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  //: IN g3 (Clk) @(93,266) /sn:0 /w:[ 0 ]
  myAND2 g2 (.b(R), .a(Clk), .out(w0));   //: @(207, 321) /sz:(89, 49) /sn:0 /p:[ Li0>1 Li1>5 Ro0<0 ]
  myAND2 g1 (.b(Clk), .a(S), .out(w2));   //: @(211, 152) /sz:(85, 47) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  //: IN g6 (R) @(83,359) /sn:0 /w:[ 0 ]
  //: OUT g7 (Y) @(580,275) /sn:0 /w:[ 0 ]
  //: IN g5 (S) @(89,159) /sn:0 /w:[ 0 ]
  //: OUT g0 (Y_n) @(553,322) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin MyINV
module MyINV(out, in);
//: interface  /sz:(98, 111) /bd:[ Li0>in(57/111) Ro0<out(56/111) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in;    //: /sn:0 {0}(223,195)(264,195){1}
//: {2}(266,193)(266,141)(275,141){3}
//: {4}(266,197)(266,227)(275,227){5}
supply1 w0;    //: /sn:0 {0}(289,87)(289,133){1}
supply0 w1;    //: /sn:0 {0}(289,272)(289,236){1}
output out;    //: /sn:0 {0}(289,219)(289,194){1}
//: {2}(291,192)(345,192){3}
//: {4}(289,190)(289,150){5}
//: enddecls

  _GGPMOS #(2, 1) g4 (.Z(out), .S(w0), .G(in));   //: @(283,141) /sn:0 /w:[ 5 1 3 ]
  //: GROUND g3 (w1) @(289,278) /sn:0 /w:[ 0 ]
  //: VDD g2 (w0) @(300,87) /sn:0 /w:[ 0 ]
  //: OUT g1 (out) @(342,192) /sn:0 /w:[ 3 ]
  //: joint g6 (in) @(266, 195) /w:[ -1 2 1 4 ]
  //: joint g7 (out) @(289, 192) /w:[ 2 4 -1 1 ]
  _GGNMOS #(2, 1) g5 (.Z(out), .S(w1), .G(in));   //: @(283,227) /sn:0 /w:[ 0 1 5 ]
  //: IN g0 (in) @(221,195) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin ControlUnit
module ControlUnit(n_clk, control, enable, clk);
//: interface  /sz:(102, 98) /bd:[ Ri0>enable(74/98) Ri1>clk(21/98) Lo0<n_clk[1:0](80/98) Lo1<control[3:0](20/98) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input enable;    //: /sn:0 {0}(794,219)(794,152){1}
//: {2}(796,150)(880,150){3}
//: {4}(792,150)(663,150)(663,217){5}
output [3:0] control;    //: /sn:0 {0}(#:910,61)(991,61){1}
output [1:0] n_clk;    //: /sn:0 {0}(186,321)(#:186,377){1}
input clk;    //: /sn:0 {0}(560,543)(560,506)(845,506)(845,417){1}
//: {2}(847,415)(906,415){3}
//: {4}(845,413)(845,319)(556,319)(556,376){5}
wire w6;    //: /sn:0 {0}(609,606)(773,606)(773,286){1}
wire w4;    //: /sn:0 {0}(605,439)(641,439)(641,284){1}
wire w0;    //: /sn:0 {0}(327,291)(327,187){1}
//: {2}(329,185)(615,185)(615,217){3}
//: {4}(327,183)(327,155)(299,155)(299,148)(370,148)(370,76)(904,76){5}
//: {6}(325,185)(281,185)(281,206)(100,206)(100,189){7}
wire w3;    //: /sn:0 {0}(509,563)(93,563)(93,281)(219,281)(219,66)(904,66){1}
wire w1;    //: /sn:0 {0}(904,46)(33,46)(33,605)(179,605){1}
//: {2}(183,605)(309,605){3}
//: {4}(313,605)(508,605){5}
//: {6}(311,603)(311,350){7}
//: {8}(181,603)(181,383){9}
wire w8;    //: /sn:0 {0}(191,383)(191,438)(450,438){1}
//: {2}(454,438)(504,438){3}
//: {4}(452,436)(452,382)(400,382){5}
//: {6}(398,380)(398,124)(746,124)(746,219){7}
//: {8}(396,382)(348,382)(348,350){9}
wire w2;    //: /sn:0 {0}(490,390)(505,390){1}
wire w9;    //: /sn:0 {0}(100,126)(100,90)(202,90)(202,56)(904,56){1}
//: enddecls

  //: comment g4 @(703,103) /sn:0
  //: /line:"S1_next"
  //: /end
  //: comment g8 @(572,165) /sn:0
  //: /line:"S0_next"
  //: /end
  //: frame g3 @(470,512) /sn:0 /wi:182 /ht:139 /tx:"S1"
  //: OUT g16 (n_clk) @(186,324) /sn:0 /R:1 /w:[ 0 ]
  assign n_clk = {w1, w8}; //: CONCAT g17  @(186,378) /sn:0 /R:1 /w:[ 1 9 0 ] /dr:0 /tp:0 /drp:1
  MyINV g26 (.in(w0), .out(w9));   //: @(68, 128) /sz:(64, 61) /R:1 /sn:0 /p:[ Bi0>7 To0<0 ]
  myFFDet g2 (.Clk(clk), .D(w6), .Y_n(w3), .Y(w1));   //: @(510, 544) /sz:(99, 80) /R:2 /sn:0 /p:[ Ti0>0 Ri0>0 Lo0<0 Lo1<5 ]
  //: comment g24 @(303,132) /sn:0
  //: /line:"d = DEMUX2"
  //: /end
  //: frame g1 @(477,348) /sn:0 /wi:182 /ht:138 /tx:"S0"
  //: joint g18 (w8) @(452, 438) /w:[ 2 4 1 -1 ]
  myAND2 g10 (.a(w8), .b(enable), .out(w6));   //: @(735, 220) /sz:(78, 65) /R:3 /sn:0 /p:[ Ti0>7 Ti1>0 Bo0<1 ]
  myNOR2 g6 (.a(w1), .b(w8), .out(w0));   //: @(299, 293) /sz:(67, 57) /R:1 /sn:0 /p:[ Bi0>7 Bi1>9 To0<0 ]
  myAND2 g9 (.a(w0), .b(enable), .out(w4));   //: @(604, 218) /sz:(77, 65) /R:3 /sn:0 /p:[ Ti0>3 Ti1>5 Bo0<1 ]
  //: joint g7 (w8) @(398, 382) /w:[ 5 6 8 -1 ]
  //: joint g22 (w0) @(327, 185) /w:[ 2 4 6 1 ]
  //: OUT g12 (control) @(988,61) /sn:0 /w:[ 1 ]
  //: comment g28 @(109,71) /sn:0
  //: /line:"b = MUX2, MUX3"
  //: /end
  //: joint g14 (enable) @(794, 150) /w:[ 2 -1 4 1 ]
  //: IN g5 (enable) @(882,150) /sn:0 /R:2 /w:[ 3 ]
  assign control = {w1, w9, w3, w0}; //: CONCAT g11  @(909,61) /sn:0 /w:[ 0 0 1 1 5 ] /dr:0 /tp:0 /drp:1
  //: joint g19 (w1) @(311, 605) /w:[ 4 6 3 -1 ]
  //: comment g21 @(37,28) /sn:0
  //: /line:"a = MUX1"
  //: /end
  //: joint g20 (w1) @(181, 605) /w:[ 2 8 1 -1 ]
  //: joint g15 (clk) @(845, 415) /w:[ 2 4 -1 1 ]
  myFFDet g0 (.Clk(clk), .D(w4), .Y_n(w2), .Y(w8));   //: @(506, 377) /sz:(99, 80) /R:2 /sn:0 /p:[ Ti0>5 Ri0>0 Lo0<1 Lo1<3 ]
  //: comment g27 @(94,259) /sn:0
  //: /line:"c = DEMUX1"
  //: /end
  //: IN g13 (clk) @(908,415) /sn:0 /R:2 /w:[ 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin myPrParziale8
module myPrParziale8(out, m, M);
//: interface  /sz:(149, 125) /bd:[ Li0>M[7:0](25/125) Li1>m(97/125) Ro0<out[7:0](62/125) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] M;    //: /sn:0 {0}(#:211,704)(211,695){1}
//: {2}(211,694)(211,610){3}
//: {4}(211,609)(211,512){5}
//: {6}(211,511)(211,419){7}
//: {8}(211,418)(211,301){9}
//: {10}(211,300)(211,211){11}
//: {12}(211,210)(211,160){13}
//: {14}(211,159)(211,85){15}
//: {16}(211,84)(211,38)(#:45,38){17}
output [7:0] out;    //: /sn:0 {0}(#:580,328)(628,328){1}
input m;    //: /sn:0 {0}(330,637)(127,637)(127,640)(117,640){1}
//: {2}(115,638)(115,545){3}
//: {4}(117,543)(127,543)(127,538)(333,538){5}
//: {6}(115,541)(115,462){7}
//: {8}(117,460)(244,460)(244,447)(333,447){9}
//: {10}(115,458)(115,351){11}
//: {12}(117,349)(127,349)(127,350)(334,350){13}
//: {14}(115,347)(115,271){15}
//: {16}(117,269)(271,269)(271,254)(336,254){17}
//: {18}(115,267)(115,196){19}
//: {20}(117,194)(151,194)(151,186)(281,186)(281,170)(334,170){21}
//: {22}(115,192)(115,118){23}
//: {24}(117,116)(269,116)(269,78)(336,78){25}
//: {26}(115,114)(115,75)(47,75){27}
//: {28}(115,642)(115,735)(329,735){29}
wire w16;    //: /sn:0 {0}(333,502)(229,502)(229,512)(215,512){1}
wire w13;    //: /sn:0 {0}(333,411)(231,411)(231,419)(215,419){1}
wire w7;    //: /sn:0 {0}(336,218)(253,218)(253,211)(215,211){1}
wire w4;    //: /sn:0 {0}(334,134)(228,134)(228,160)(215,160){1}
wire w22;    //: /sn:0 {0}(329,699)(204,699)(204,695)(206,695){1}
wire w0;    //: /sn:0 {0}(336,42)(227,42)(227,85)(215,85){1}
wire w20;    //: /sn:0 {0}(574,353)(507,353)(507,621)(413,621){1}
wire w19;    //: /sn:0 {0}(330,601)(234,601)(234,610)(215,610){1}
wire w23;    //: /sn:0 {0}(574,363)(525,363)(525,719)(412,719){1}
wire w10;    //: /sn:0 {0}(334,314)(204,314)(204,301)(206,301){1}
wire w8;    //: /sn:0 {0}(574,313)(455,313)(455,238)(419,238){1}
wire w17;    //: /sn:0 {0}(574,343)(488,343)(488,522)(416,522){1}
wire w14;    //: /sn:0 {0}(574,333)(468,333)(468,431)(416,431){1}
wire w11;    //: /sn:0 {0}(574,323)(456,323)(456,334)(417,334){1}
wire w2;    //: /sn:0 {0}(419,63)(549,63)(549,293)(574,293){1}
wire w5;    //: /sn:0 {0}(574,303)(501,303)(501,154)(417,154){1}
//: enddecls

  myAND2 g8 (.b(m), .a(w22), .out(w23));   //: @(330, 690) /sz:(81, 59) /sn:0 /p:[ Li0>29 Li1>0 Ro0<1 ]
  myAND2 g4 (.b(m), .a(w10), .out(w11));   //: @(335, 305) /sz:(81, 59) /sn:0 /p:[ Li0>13 Li1>0 Ro0<1 ]
  assign w22 = M[7]; //: TAP g16 @(209,695) /sn:0 /R:2 /w:[ 1 1 2 ] /ss:0
  myAND2 g3 (.b(m), .a(w7), .out(w8));   //: @(337, 209) /sz:(81, 59) /sn:0 /p:[ Li0>17 Li1>0 Ro0<1 ]
  //: OUT g26 (out) @(625,328) /sn:0 /w:[ 1 ]
  //: IN g17 (m) @(45,75) /sn:0 /w:[ 27 ]
  myAND2 g2 (.b(m), .a(w4), .out(w5));   //: @(335, 125) /sz:(81, 59) /sn:0 /p:[ Li0>21 Li1>0 Ro0<1 ]
  //: joint g23 (m) @(115, 543) /w:[ 4 6 -1 3 ]
  //: joint g24 (m) @(115, 640) /w:[ 1 2 -1 28 ]
  //: IN g1 (M) @(43,38) /sn:0 /w:[ 17 ]
  //: joint g18 (m) @(115, 116) /w:[ 24 26 -1 23 ]
  assign out = {w23, w20, w17, w14, w11, w8, w5, w2}; //: CONCAT g25  @(579,328) /sn:0 /w:[ 0 0 0 0 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  assign w4 = M[1]; //: TAP g10 @(209,160) /sn:0 /R:2 /w:[ 1 13 14 ] /ss:1
  myAND2 g6 (.b(m), .a(w16), .out(w17));   //: @(334, 493) /sz:(81, 59) /sn:0 /p:[ Li0>5 Li1>0 Ro0<1 ]
  assign w0 = M[0]; //: TAP g9 @(209,85) /sn:0 /R:2 /w:[ 1 15 16 ] /ss:1
  myAND2 g7 (.b(m), .a(w19), .out(w20));   //: @(331, 592) /sz:(81, 59) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: joint g22 (m) @(115, 460) /w:[ 8 10 -1 7 ]
  assign w10 = M[3]; //: TAP g12 @(209,301) /sn:0 /R:2 /w:[ 1 9 10 ] /ss:0
  assign w16 = M[5]; //: TAP g14 @(209,512) /sn:0 /R:2 /w:[ 1 5 6 ] /ss:1
  assign w7 = M[2]; //: TAP g11 @(209,211) /sn:0 /R:2 /w:[ 1 11 12 ] /ss:1
  myAND2 g5 (.b(m), .a(w13), .out(w14));   //: @(334, 402) /sz:(81, 59) /sn:0 /p:[ Li0>9 Li1>0 Ro0<1 ]
  //: joint g21 (m) @(115, 349) /w:[ 12 14 -1 11 ]
  //: joint g19 (m) @(115, 194) /w:[ 20 22 -1 19 ]
  //: joint g20 (m) @(115, 269) /w:[ 16 18 -1 15 ]
  assign w19 = M[6]; //: TAP g15 @(209,610) /sn:0 /R:2 /w:[ 1 3 4 ] /ss:1
  myAND2 g0 (.b(m), .a(w0), .out(w2));   //: @(337, 33) /sz:(81, 59) /sn:0 /p:[ Li0>25 Li1>0 Ro0<0 ]
  assign w13 = M[4]; //: TAP g13 @(209,419) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin myADD8
module myADD8(A, Cin, S, B, Cout);
//: interface  /sz:(77, 220) /bd:[ Ti0>Cin(40/77) Li0>B[7:0](172/220) Li1>A[7:0](41/220) Bo0<Cout(39/77) Ro0<S[7:0](102/220) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] B;    //: /sn:0 {0}(#:76,29)(161,29){1}
//: {2}(162,29)(301,29){3}
//: {4}(302,29)(502,29){5}
//: {6}(503,29)(656,29){7}
//: {8}(657,29)(813,29){9}
//: {10}(814,29)(1009,29){11}
//: {12}(1010,29)(1178,29){13}
//: {14}(1179,29)(1357,29){15}
//: {16}(1358,29)(1448,29){17}
input [7:0] A;    //: /sn:0 {0}(#:78,77)(193,77){1}
//: {2}(194,77)(346,77){3}
//: {4}(347,77)(553,77){5}
//: {6}(554,77)(727,77){7}
//: {8}(728,77)(853,77){9}
//: {10}(854,77)(1062,77){11}
//: {12}(1063,77)(1248,77){13}
//: {14}(1249,77)(1398,77){15}
//: {16}(1399,77)(1438,77){17}
input Cin;    //: /sn:0 {0}(1519,78)(1519,227)(1419,227){1}
output Cout;    //: /sn:0 {0}(148,235)(69,235){1}
output [7:0] S;    //: /sn:0 {0}(163,380)(#:197,380){1}
wire w6;    //: /sn:0 {0}(203,365)(524,365)(524,270){1}
wire w13;    //: /sn:0 {0}(1221,228)(1320,228){1}
wire w16;    //: /sn:0 {0}(1249,81)(1249,129)(1200,129)(1200,199){1}
wire w7;    //: /sn:0 {0}(203,375)(685,375)(685,267){1}
wire w34;    //: /sn:0 {0}(162,33)(162,97)(164,97)(164,204){1}
wire w4;    //: /sn:0 {0}(358,270)(358,355)(203,355){1}
wire w25;    //: /sn:0 {0}(657,33)(657,39)(651,39)(651,196){1}
wire w36;    //: /sn:0 {0}(1371,264)(1371,415)(203,415){1}
wire w3;    //: /sn:0 {0}(203,345)(273,345)(273,291)(194,291)(194,271){1}
wire w0;    //: /sn:0 {0}(573,229)(633,229){1}
wire w22;    //: /sn:0 {0}(897,230)(957,230){1}
wire w20;    //: /sn:0 {0}(1063,81)(1063,106)(1035,106)(1035,201){1}
wire w30;    //: /sn:0 {0}(302,33)(302,39)(328,39)(328,201){1}
wire w29;    //: /sn:0 {0}(503,33)(503,111)(491,111)(491,197){1}
wire w18;    //: /sn:0 {0}(1056,229)(1122,229){1}
wire w19;    //: /sn:0 {0}(203,405)(1173,405)(1173,265){1}
wire w23;    //: /sn:0 {0}(203,395)(1008,395)(1008,265){1}
wire w10;    //: /sn:0 {0}(1358,33)(1358,134)(1338,134)(1338,198){1}
wire w24;    //: /sn:0 {0}(854,81)(854,89)(876,89)(876,198){1}
wire w21;    //: /sn:0 {0}(814,33)(814,41)(816,41)(816,198){1}
wire w1;    //: /sn:0 {0}(405,231)(473,231){1}
wire w32;    //: /sn:0 {0}(554,81)(554,137)(551,137)(551,197){1}
wire w8;    //: /sn:0 {0}(849,272)(849,385)(203,385){1}
wire w17;    //: /sn:0 {0}(1010,33)(1010,110)(975,110)(975,201){1}
wire w33;    //: /sn:0 {0}(347,81)(347,87)(385,87)(385,201){1}
wire w28;    //: /sn:0 {0}(728,81)(728,146)(713,146)(713,196){1}
wire w2;    //: /sn:0 {0}(240,233)(312,233){1}
wire w11;    //: /sn:0 {0}(1399,81)(1399,96)(1398,96)(1398,198){1}
wire w15;    //: /sn:0 {0}(1179,33)(1179,136)(1140,136)(1140,199){1}
wire w38;    //: /sn:0 {0}(194,81)(194,134)(220,134)(220,204){1}
wire w26;    //: /sn:0 {0}(798,232)(735,232){1}
//: enddecls

  myFA g8 (.B(w29), .A(w32), .Cin(w0), .Cout(w1), .S(w6));   //: @(474, 198) /sz:(98, 71) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  myFA g4 (.B(w15), .A(w16), .Cin(w13), .Cout(w18), .S(w19));   //: @(1123, 200) /sz:(97, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  assign w28 = A[4]; //: TAP g16 @(728,75) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  myFA g3 (.B(w10), .A(w11), .Cin(Cin), .Cout(w13), .S(w36));   //: @(1321, 199) /sz:(97, 64) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  assign w21 = B[3]; //: TAP g26 @(814,27) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  assign w24 = A[3]; //: TAP g17 @(854,75) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  //: IN g2 (A) @(76,77) /sn:0 /w:[ 0 ]
  assign w30 = B[6]; //: TAP g23 @(302,27) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w29 = B[5]; //: TAP g24 @(503,27) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: IN g1 (Cin) @(1519,76) /sn:0 /R:3 /w:[ 0 ]
  assign w10 = B[0]; //: TAP g29 @(1358,27) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign w20 = A[2]; //: TAP g18 @(1063,75) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  assign w25 = B[4]; //: TAP g25 @(657,27) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  myFA g10 (.B(w34), .A(w38), .Cin(w2), .Cout(Cout), .S(w3));   //: @(149, 205) /sz:(90, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<1 ]
  myFA g6 (.B(w21), .A(w24), .Cin(w22), .Cout(w26), .S(w8));   //: @(799, 199) /sz:(97, 72) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  myFA g9 (.B(w30), .A(w33), .Cin(w1), .Cout(w2), .S(w4));   //: @(313, 202) /sz:(91, 67) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  myFA g7 (.B(w25), .A(w28), .Cin(w26), .Cout(w0), .S(w7));   //: @(634, 197) /sz:(100, 69) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  assign w34 = B[7]; //: TAP g22 @(162,27) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: OUT g12 (S) @(166,380) /sn:0 /R:2 /w:[ 0 ]
  assign w15 = B[1]; //: TAP g28 @(1179,27) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  assign w33 = A[6]; //: TAP g14 @(347,75) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w38 = A[7]; //: TAP g11 @(194,75) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  myFA g5 (.B(w17), .A(w20), .Cin(w18), .Cout(w22), .S(w23));   //: @(958, 202) /sz:(97, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: IN g21 (B) @(74,29) /sn:0 /w:[ 0 ]
  assign w16 = A[1]; //: TAP g19 @(1249,75) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  assign w11 = A[0]; //: TAP g20 @(1399,75) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  assign w32 = A[5]; //: TAP g15 @(554,75) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: OUT g0 (Cout) @(72,235) /sn:0 /R:2 /w:[ 1 ]
  assign w17 = B[2]; //: TAP g27 @(1010,27) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  assign S = {w3, w4, w6, w7, w8, w23, w19, w36}; //: CONCAT g13  @(198,380) /sn:0 /R:2 /w:[ 1 0 1 0 0 1 0 0 1 ] /dr:0 /tp:0 /drp:1

endmodule
//: /netlistEnd

//: /netlistBegin myHA
module myHA(out, b, a, cout);
//: interface  /sz:(85, 110) /bd:[ Li0>b(87/110) Li1>a(20/110) Ri0>out(50/110) Bo0<cout(43/85) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(271,193)(205,193)(205,328){1}
//: {2}(207,330)(275,330){3}
//: {4}(203,330)(150,330){5}
output out;    //: /sn:0 {0}(358,163)(464,163){1}
output cout;    //: /sn:0 {0}(379,307)(455,307){1}
input a;    //: /sn:0 {0}(275,280)(185,280)(185,131){1}
//: {2}(187,129)(271,129){3}
//: {4}(185,127)(185,91)(137,91){5}
//: enddecls

  //: OUT g4 (out) @(461,163) /sn:0 /w:[ 1 ]
  //: IN g3 (b) @(148,330) /sn:0 /w:[ 5 ]
  //: IN g2 (a) @(135,91) /sn:0 /w:[ 5 ]
  myAND2 g1 (.a(a), .b(b), .out(cout));   //: @(276, 267) /sz:(102, 81) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  //: joint g6 (a) @(185, 129) /w:[ 2 4 -1 1 ]
  //: joint g7 (b) @(205, 330) /w:[ 2 1 4 -1 ]
  //: OUT g5 (cout) @(452,307) /sn:0 /w:[ 1 ]
  myXOR g0 (.A(a), .B(b), .out(out));   //: @(272, 109) /sz:(85, 111) /sn:0 /p:[ Li0>3 Li1>0 Ro0<0 ]

endmodule
//: /netlistEnd

