//: version "2.1"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "MUX2.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] w19;    //: /sn:0 {0}(359,102)(266,102)(#:266,94){1}
reg [3:0] w21;    //: /sn:0 {0}(#:265,143)(265,153)(359,153){1}
reg w1;    //: /sn:0 {0}(409,40)(409,79){1}
reg w5;    //: /sn:0 {0}(412,237)(412,178){1}
wire [15:0] S;    //: /sn:0 {0}(#:550,116)(550,124)(459,124){1}
//: enddecls

  //: DIP g3 (w19) @(266,84) /sn:0 /w:[ 1 ] /st:2 /dn:0
  //: SWITCH g16 (w5) @(412,251) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:0
  //: SWITCH g18 (w1) @(409,27) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:0
  //: DIP g9 (w21) @(265,133) /sn:0 /w:[ 0 ] /st:3 /dn:0
  //: LED g20 (S) @(550,109) /sn:0 /w:[ 0 ] /type:3
  QUADRATO g0 (.Clk(w1), .B(w21), .A(w19), .Start(w5), .S(S));   //: @(360, 80) /sz:(98, 97) /sn:0 /p:[ Ti0>1 Li0>1 Li1>0 Bi0>1 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin EXOR2
module EXOR2(b, out, a);
//: interface  /sz:(45, 43) /bd:[ Li0>a(10/43) Li1>b(30/43) Ro0<out(21/43) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(38,192)(52,192){1}
//: {2}(56,192)(92,192){3}
//: {4}(54,190)(54,130)(172,130)(172,107)(203,107){5}
output out;    //: /sn:0 {0}(330,134)(370,134){1}
input a;    //: /sn:0 {0}(206,171)(173,171)(173,151)(68,151)(68,90){1}
//: {2}(70,88)(93,88){3}
//: {4}(66,88)(40,88){5}
wire w6;    //: /sn:0 {0}(245,95)(273,95)(273,126)(288,126){1}
wire w3;    //: /sn:0 {0}(134,191)(206,191){1}
wire w1;    //: /sn:0 {0}(135,87)(203,87){1}
wire w9;    //: /sn:0 {0}(248,179)(273,179)(273,146)(288,146){1}
//: enddecls

  //: joint g8 (a) @(68, 88) /w:[ 2 -1 4 1 ]
  NAND2 g4 (.in2(b), .in1(w1), .out(w6));   //: @(204, 77) /sz:(40, 40) /sn:0 /p:[ Li0>5 Li1>1 Ro0<0 ]
  INV1 g3 (.in(b), .out(w3));   //: @(93, 171) /sz:(40, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  INV1 g2 (.in(a), .out(w1));   //: @(94, 67) /sz:(40, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: IN g1 (b) @(36,192) /sn:0 /w:[ 0 ]
  //: joint g6 (b) @(54, 192) /w:[ 2 4 1 -1 ]
  //: OUT g9 (out) @(367,134) /sn:0 /w:[ 1 ]
  NAND2 g7 (.in2(w9), .in1(w6), .out(out));   //: @(289, 116) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  NAND2 g5 (.in2(w3), .in1(a), .out(w9));   //: @(207, 161) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  //: IN g0 (a) @(38,88) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin QUADRATO
module QUADRATO(Clk, A, S, B, Start);
//: interface  /sz:(98, 97) /bd:[ Ti0>Clk(49/98) Li0>B[7:0](73/97) Li1>A[7:0](22/97) Bi0>Start(52/98) Ro0<S[15:0](44/97) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input Start;    //: /sn:0 {0}(181,6)(181,-51){1}
input [3:0] B;    //: /sn:0 {0}(#:403,-147)(403,-111){1}
supply0 [7:0] w25;    //: /sn:0 {0}(#:348,468)(348,501)(#:375,501){1}
input [3:0] A;    //: /sn:0 {0}(287,-116)(#:287,-145){1}
supply0 [3:0] w0;    //: /sn:0 {0}(#:326,15)(312,15)(#:312,33){1}
input Clk;    //: /sn:0 {0}(312,382)(139,382)(139,31){1}
//: {2}(141,29)(154,29){3}
//: {4}(139,27)(139,-15){5}
//: {6}(141,-17)(444,-17)(444,-73)(429,-73){7}
//: {8}(139,-19)(139,-27){9}
//: {10}(141,-29)(325,-29)(325,-78)(313,-78){11}
//: {12}(139,-31)(139,-49){13}
supply0 [3:0] w14;    //: /sn:0 {0}(#:447,17)(428,17)(#:428,33){1}
output [15:0] S;    //: /sn:0 {0}(#:343,415)(343,430){1}
//: {2}(345,432)(549,432)(549,430)(#:553,430){3}
//: {4}(343,434)(#:343,462){5}
wire [7:0] w16;    //: /sn:0 {0}(#:292,39)(#:292,97){1}
wire w13;    //: /sn:0 {0}(418,1)(418,33){1}
wire w6;    //: /sn:0 {0}(272,-1)(272,33){1}
wire w7;    //: /sn:0 {0}(282,-1)(282,33){1}
wire [7:0] w4;    //: /sn:0 {0}(#:280,139)(280,178)(331,178)(#:331,215){1}
wire [15:0] w3;    //: /sn:0 {0}(343,349)(#:343,280){1}
wire [7:0] w20;    //: /sn:0 {0}(#:408,39)(#:408,98){1}
wire w12;    //: /sn:0 {0}(408,1)(408,33){1}
wire [3:0] w19;    //: /sn:0 {0}(403,-34)(#:403,-5){1}
wire w10;    //: /sn:0 {0}(388,1)(388,33){1}
wire w1;    //: /sn:0 {0}(305,117)(343,117)(343,198){1}
//: {2}(345,200)(456,200)(456,118)(421,118){3}
//: {4}(341,200)(188,200)(188,60){5}
wire w8;    //: /sn:0 {0}(292,-1)(292,33){1}
wire [7:0] w17;    //: /sn:0 {0}(#:338,468)(338,526){1}
//: {2}(340,528)(479,528)(#:479,68)(382,68)(#:382,98){3}
//: {4}(336,528)(213,528)(213,66)(266,66)(#:266,97){5}
wire [7:0] w2;    //: /sn:0 {0}(#:361,215)(361,178)(396,178)(#:396,140){1}
wire w11;    //: /sn:0 {0}(398,1)(398,33){1}
wire [3:0] w5;    //: /sn:0 {0}(287,-39)(#:287,-7){1}
wire w9;    //: /sn:0 {0}(302,-1)(302,33){1}
//: enddecls

  assign w20 = {w14, w13, w12, w11, w10}; //: CONCAT g8  @(408,38) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  assign {w9, w8, w7, w6} = w5; //: CONCAT g4  @(287,-6) /sn:0 /R:1 /w:[ 0 0 0 0 1 ] /dr:1 /tp:0 /drp:0
  //: IN g16 (Clk) @(139,-51) /sn:0 /R:3 /w:[ 13 ]
  //: IN g3 (A) @(287,-147) /sn:0 /R:3 /w:[ 1 ]
  //: OUT g17 (S) @(550,430) /sn:0 /w:[ 3 ]
  //: GROUND g2 (w0) @(332,15) /sn:0 /R:1 /w:[ 0 ]
  //: joint g23 (Clk) @(139, -17) /w:[ 6 8 -1 5 ]
  CU g24 (.in(Start), .Clk(Clk), .out(w1));   //: @(155, 7) /sz:(63, 52) /sn:0 /p:[ Ti0>0 Li0>3 Bo0<5 ]
  assign w16 = {w0, w9, w8, w7, w6}; //: CONCAT g1  @(292,38) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  REG4 g18 (.in(A), .Clk(Clk), .out(w5));   //: @(260, -115) /sz:(52, 75) /R:3 /sn:0 /p:[ Ti0>0 Ri0>11 Bo0<0 ]
  //: joint g25 (w1) @(343, 200) /w:[ 2 1 4 -1 ]
  MUX8 g10 (.b(w17), .a(w16), .C(w1), .out(w4));   //: @(254, 98) /sz:(50, 40) /R:3 /sn:0 /p:[ Ti0>5 Ti1>1 Ri0>0 Bo0<0 ]
  //: joint g6 (w17) @(338, 528) /w:[ 2 1 4 -1 ]
  //: IN g9 (B) @(403,-149) /sn:0 /R:3 /w:[ 0 ]
  //: GROUND g7 (w14) @(453,17) /sn:0 /R:1 /w:[ 0 ]
  //: joint g22 (Clk) @(139, -29) /w:[ 10 12 -1 9 ]
  REG16 g12 (.in(w3), .clk(Clk), .out(S));   //: @(314, 350) /sz:(59, 64) /R:3 /sn:0 /p:[ Ti0>0 Li0>0 Bo0<0 ]
  //: GROUND g14 (w25) @(381,501) /sn:0 /R:1 /w:[ 1 ]
  MUX8 g11 (.b(w17), .a(w20), .C(w1), .out(w2));   //: @(370, 99) /sz:(50, 40) /R:3 /sn:0 /p:[ Ti0>3 Ti1>1 Ri0>3 Bo0<1 ]
  assign {w13, w12, w11, w10} = w19; //: CONCAT g5  @(403,-4) /sn:0 /R:1 /w:[ 0 0 0 0 1 ] /dr:1 /tp:0 /drp:0
  REG4 g21 (.in(B), .Clk(Clk), .out(w19));   //: @(376, -110) /sz:(52, 75) /R:3 /sn:0 /p:[ Ti0>1 Ri0>7 Bo0<0 ]
  //: joint g19 (Clk) @(139, 29) /w:[ 2 4 -1 1 ]
  //: IN g20 (Start) @(181,-53) /sn:0 /R:3 /w:[ 1 ]
  MUL8 g0 (.a(w2), .b(w4), .out(w3));   //: @(313, 216) /sz:(62, 63) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<1 ]
  //: joint g15 (S) @(343, 432) /w:[ 2 1 -1 4 ]
  assign {w25, w17} = S; //: CONCAT g13  @(343,463) /sn:0 /R:1 /w:[ 0 0 5 ] /dr:1 /tp:1 /drp:0

endmodule
//: /netlistEnd

//: /netlistBegin FFSR
module FFSR(S, Y, clk, R);
//: interface  /sz:(40, 40) /bd:[ Li0>R(28/40) Li1>S(7/40) Bi0>clk(17/40) Ro0<Y(18/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input R;    //: /sn:0 {0}(300,174)(215,174){1}
input clk;    //: /sn:0 {0}(300,194)(267,194){1}
//: {2}(265,192)(265,127)(301,127){3}
//: {4}(265,196)(265,238){5}
supply0 w2;    //: /sn:0 {0}(479,154)(507,154){1}
input S;    //: /sn:0 {0}(214,107)(301,107){1}
output Y;    //: /sn:0 {0}(479,175)(514,175){1}
wire w0;    //: /sn:0 {0}(342,183)(381,183)(381,175)(396,175){1}
wire w1;    //: /sn:0 {0}(343,116)(381,116)(381,151)(396,151){1}
//: enddecls

  //: IN g4 (S) @(212,107) /sn:0 /w:[ 0 ]
  //: GROUND g8 (w2) @(513,154) /sn:0 /R:1 /w:[ 1 ]
  AND2 g3 (.in2(clk), .in1(S), .out(w1));   //: @(302, 97) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  AND2 g2 (.in2(clk), .in1(R), .out(w0));   //: @(301, 164) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: OUT g1 (Y) @(511,175) /sn:0 /w:[ 1 ]
  //: IN g6 (clk) @(265,240) /sn:0 /R:1 /w:[ 5 ]
  //: joint g7 (clk) @(265, 194) /w:[ 1 2 -1 4 ]
  //: IN g5 (R) @(213,174) /sn:0 /w:[ 1 ]
  LATCHSR g0 (.s(w1), .r(w0), .Y1(w2), .Y(Y));   //: @(397, 144) /sz:(81, 47) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA4
module FA4(s, b, cin, cout, a);
//: interface  /sz:(40, 40) /bd:[ Ti0>b[3:0](28/40) Ti1>a[3:0](10/40) Ri0>cin(19/40) Lo0<cout(19/40) Bo0<s[3:0](17/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:761,200)(657,200){1}
//: {2}(656,200)(524,200){3}
//: {4}(523,200)(388,200){5}
//: {6}(387,200)(247,200){7}
//: {8}(246,200)(#:236,200){9}
input cin;    //: /sn:0 {0}(707,285)(767,285){1}
output cout;    //: /sn:0 {0}(228,281)(185,281){1}
output [3:0] s;    //: /sn:0 {0}(468,451)(#:468,420){1}
input [3:0] a;    //: /sn:0 {0}(#:757,158)(688,158){1}
//: {2}(687,158)(555,158){3}
//: {4}(554,158)(419,158){5}
//: {6}(418,158)(278,158){7}
//: {8}(277,158)(#:269,158){9}
wire w6;    //: /sn:0 {0}(419,249)(419,162){1}
wire w16;    //: /sn:0 {0}(688,251)(688,162){1}
wire w13;    //: /sn:0 {0}(463,414)(463,387)(400,387)(400,313){1}
wire w7;    //: /sn:0 {0}(369,282)(297,282){1}
wire w4;    //: /sn:0 {0}(259,312)(259,396)(453,396)(453,414){1}
wire w0;    //: /sn:0 {0}(278,248)(278,162){1}
wire w3;    //: /sn:0 {0}(555,162)(555,250){1}
wire w19;    //: /sn:0 {0}(483,414)(483,396)(669,396)(669,315){1}
wire w1;    //: /sn:0 {0}(247,248)(247,204){1}
wire w8;    //: /sn:0 {0}(438,283)(505,283){1}
wire w17;    //: /sn:0 {0}(536,314)(536,387)(473,387)(473,414){1}
wire w2;    //: /sn:0 {0}(524,204)(524,250){1}
wire w15;    //: /sn:0 {0}(657,251)(657,204){1}
wire w5;    //: /sn:0 {0}(388,249)(388,204){1}
wire w9;    //: /sn:0 {0}(638,284)(574,284){1}
//: enddecls

  assign w3 = a[1]; //: TAP g8 @(555,156) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  FA2 g4 (.b(w6), .a(w5), .cin(w8), .cout(w7), .s(w13));   //: @(370, 250) /sz:(67, 62) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  assign w0 = a[3]; //: TAP g3 @(278,156) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  assign s = {w4, w13, w17, w19}; //: CONCAT g16  @(468,419) /sn:0 /R:3 /w:[ 1 1 0 1 0 ] /dr:1 /tp:0 /drp:1
  //: OUT g17 (s) @(468,448) /sn:0 /R:3 /w:[ 0 ]
  FA2 g2 (.b(w0), .a(w1), .cin(w7), .cout(cout), .s(w4));   //: @(229, 249) /sz:(67, 62) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  //: IN g1 (b) @(763,200) /sn:0 /R:2 /w:[ 0 ]
  assign w1 = b[3]; //: TAP g10 @(247,198) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  FA2 g6 (.a(w15), .b(w16), .cin(cin), .cout(w9), .s(w19));   //: @(639, 252) /sz:(67, 62) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  assign w6 = a[2]; //: TAP g7 @(419,156) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  assign w16 = a[0]; //: TAP g9 @(688,156) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  assign w2 = b[1]; //: TAP g12 @(524,198) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  assign w5 = b[2]; //: TAP g11 @(388,198) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: IN g14 (cin) @(769,285) /sn:0 /R:2 /w:[ 1 ]
  FA2 g5 (.b(w3), .a(w2), .cin(w9), .cout(w8), .s(w17));   //: @(506, 251) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  //: OUT g15 (cout) @(188,281) /sn:0 /R:2 /w:[ 1 ]
  //: IN g0 (a) @(759,158) /sn:0 /R:2 /w:[ 0 ]
  assign w15 = b[0]; //: TAP g13 @(657,198) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin CU
module CU(out, Clk, in);
//: interface  /sz:(63, 52) /bd:[ Ti0>in(26/63) Li0>Clk(22/52) Bo0<out(33/63) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input in;    //: /sn:0 {0}(499,634)(499,519){1}
//: {2}(499,515)(499,454)(457,454){3}
//: {4}(497,517)(458,517){5}
input Clk;    //: /sn:0 {0}(627,473)(627,463)(588,463){1}
//: {2}(586,461)(586,396)(629,396)(629,410){3}
//: {4}(586,465)(586,637){5}
output out;    //: /sn:0 {0}(300,175)(221,175){1}
//: {2}(219,173)(219,67)(730,67){3}
//: {4}(734,67)(786,67){5}
//: {6}(732,69)(732,495)(646,495){7}
//: {8}(219,177)(219,445)(310,445){9}
wire w6;    //: /sn:0 {0}(461,182)(526,182)(526,155)(541,155){1}
wire w7;    //: /sn:0 {0}(462,109)(526,109)(526,135)(541,135){1}
wire w0;    //: /sn:0 {0}(583,143)(690,143)(690,432)(648,432){1}
wire w12;    //: /sn:0 {0}(419,194)(199,194){1}
//: {2}(197,192)(197,102)(301,102){3}
//: {4}(197,196)(197,508)(309,508){5}
wire w10;    //: /sn:0 {0}(343,101)(420,101){1}
wire w21;    //: /sn:0 {0}(352,444)(415,444){1}
wire w24;    //: /sn:0 {0}(351,507)(416,507){1}
wire w2;    //: /sn:0 {0}(458,495)(604,495){1}
wire w5;    //: /sn:0 {0}(457,432)(606,432){1}
wire w9;    //: /sn:0 {0}(420,121)(381,121)(381,172){1}
//: {2}(383,174)(419,174){3}
//: {4}(379,174)(342,174){5}
//: enddecls

  NAND2 g4 (.in1(w9), .in2(w12), .out(w6));   //: @(420, 164) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>0 Ro0<0 ]
  NOR2 g8 (.in2(w2), .in1(in), .out(w24));   //: @(417, 485) /sz:(40, 40) /R:2 /sn:0 /p:[ Ri0>0 Ri1>5 Lo0<1 ]
  NAND2 g3 (.in1(w10), .in2(w9), .out(w7));   //: @(421, 91) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  //: joint g16 (out) @(219, 175) /w:[ 1 2 -1 8 ]
  //: joint g17 (out) @(732, 67) /w:[ 4 -1 3 6 ]
  NAND2 g2 (.in1(w7), .in2(w6), .out(w0));   //: @(542, 125) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  FFD g1 (.Clk(Clk), .D(out), .Y(w2));   //: @(605, 474) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>0 Ri0>7 Lo0<1 ]
  //: OUT g18 (out) @(783,67) /sn:0 /w:[ 5 ]
  INV1 g10 (.in(w24), .out(w12));   //: @(310, 488) /sz:(40, 40) /R:2 /sn:0 /p:[ Ri0>0 Lo0<5 ]
  INV1 g6 (.in(out), .out(w9));   //: @(301, 154) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<5 ]
  NOR2 g7 (.in2(w5), .in1(in), .out(w21));   //: @(416, 422) /sz:(40, 40) /R:2 /sn:0 /p:[ Ri0>0 Ri1>3 Lo0<1 ]
  INV1 g9 (.in(w21), .out(out));   //: @(311, 425) /sz:(40, 40) /R:2 /sn:0 /p:[ Ri0>0 Lo0<9 ]
  //: joint g12 (w9) @(381, 174) /w:[ 2 1 4 -1 ]
  //: IN g11 (Clk) @(586,639) /sn:0 /R:1 /w:[ 5 ]
  INV1 g5 (.in(w12), .out(w10));   //: @(302, 81) /sz:(40, 40) /sn:0 /p:[ Li0>3 Ro0<0 ]
  //: joint g14 (w12) @(197, 194) /w:[ 1 2 -1 4 ]
  //: joint g19 (in) @(499, 517) /w:[ -1 2 4 1 ]
  //: joint g15 (Clk) @(586, 463) /w:[ 1 2 -1 4 ]
  FFD g0 (.Clk(Clk), .D(w0), .Y(w5));   //: @(607, 411) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>3 Ri0>1 Lo0<1 ]
  //: IN g13 (in) @(499,636) /sn:0 /R:1 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin LATCHSR
module LATCHSR(Y1, r, s, Y);
//: interface  /sz:(81, 47) /bd:[ Li0>s(7/47) Li1>r(31/47) Ro0<Y1(10/47) Ro1<Y(31/47) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input r;    //: /sn:0 {0}(253,213)(197,213){1}
input s;    //: /sn:0 {0}(255,113)(199,113){1}
output Y1;    //: /sn:0 {0}(297,123)(333,123){1}
//: {2}(337,123)(386,123){3}
//: {4}(335,125)(335,167)(243,167)(243,191)(253,191){5}
output Y;    //: /sn:0 {0}(255,135)(246,135)(246,157)(319,157)(319,199){1}
//: {2}(321,201)(381,201){3}
//: {4}(317,201)(295,201){5}
//: enddecls

  //: OUT g4 (Y1) @(383,123) /sn:0 /w:[ 3 ]
  //: IN g3 (r) @(195,213) /sn:0 /w:[ 1 ]
  //: IN g2 (s) @(197,113) /sn:0 /w:[ 1 ]
  NOR2 g1 (.in2(r), .in1(Y1), .out(Y));   //: @(254, 183) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>5 Ro0<5 ]
  //: joint g6 (Y) @(319, 201) /w:[ 2 1 4 -1 ]
  //: joint g7 (Y1) @(335, 123) /w:[ 2 -1 1 4 ]
  //: OUT g5 (Y) @(378,201) /sn:0 /w:[ 3 ]
  NOR2 g0 (.in2(Y), .in1(s), .out(Y1));   //: @(256, 105) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA2
module FA2(cout, a, b, cin, s);
//: interface  /sz:(67, 62) /bd:[ Ti0>b(49/67) Ti1>a(18/67) Ri0>cin(33/62) Lo0<cout(32/62) Bo0<s(30/67) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(71,296)(146,296){1}
//: {2}(150,296)(228,296){3}
//: {4}(148,294)(148,147)(227,147){5}
input cin;    //: /sn:0 {0}(348,337)(344,337)(344,230){1}
//: {2}(344,226)(344,192)(357,192){3}
//: {4}(342,228)(72,228){5}
output cout;    //: /sn:0 {0}(491,292)(533,292){1}
output s;    //: /sn:0 {0}(440,183)(404,183){1}
input a;    //: /sn:0 {0}(228,276)(116,276)(116,129){1}
//: {2}(118,127)(227,127){3}
//: {4}(114,127)(64,127){5}
wire w10;    //: /sn:0 {0}(390,345)(422,345)(422,304)(449,304){1}
wire w1;    //: /sn:0 {0}(348,357)(306,357)(306,140){1}
//: {2}(308,138)(342,138)(342,172)(357,172){3}
//: {4}(304,138)(274,138){5}
wire w8;    //: /sn:0 {0}(270,284)(449,284){1}
//: enddecls

  NAND2 g4 (.in1(w8), .in2(w10), .out(cout));   //: @(450, 274) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: OUT g8 (cout) @(530,292) /sn:0 /w:[ 1 ]
  //: IN g3 (a) @(62,127) /sn:0 /w:[ 5 ]
  EXOR2 g2 (.b(cin), .a(w1), .out(s));   //: @(358, 162) /sz:(45, 43) /sn:0 /p:[ Li0>3 Li1>3 Ro0<1 ]
  NAND2 g1 (.in1(a), .in2(b), .out(w8));   //: @(229, 266) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  //: joint g10 (w1) @(306, 138) /w:[ 2 -1 4 1 ]
  //: IN g6 (b) @(69,296) /sn:0 /w:[ 0 ]
  //: joint g9 (cin) @(344, 228) /w:[ -1 2 4 1 ]
  //: IN g7 (cin) @(70,228) /sn:0 /w:[ 5 ]
  //: joint g11 (a) @(116, 127) /w:[ 2 -1 4 1 ]
  EXOR2 g14 (.b(b), .a(a), .out(w1));   //: @(228, 117) /sz:(45, 43) /sn:0 /p:[ Li0>5 Li1>3 Ro0<5 ]
  NAND2 g5 (.in1(cin), .in2(w1), .out(w10));   //: @(349, 327) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: joint g0 (b) @(148, 296) /w:[ 2 4 1 -1 ]
  //: OUT g13 (s) @(437,183) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFDLS
module FFDLS(Clk, D, Y);
//: interface  /sz:(40, 40) /bd:[ Li0>D(19/40) Bi0>Clk(18/40) Ro0<Y(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(374,178)(374,148){1}
input D;    //: /sn:0 {0}(268,145)(215,145)(215,116){1}
//: {2}(217,114)(356,114){3}
//: {4}(215,112)(215,114)(194,114){5}
output Y;    //: /sn:0 {0}(398,125)(427,125){1}
wire w0;    //: /sn:0 {0}(356,135)(320,135)(320,144)(310,144){1}
//: enddecls

  //: IN g4 (Clk) @(374,180) /sn:0 /R:1 /w:[ 0 ]
  //: joint g3 (D) @(215, 114) /w:[ 2 4 -1 1 ]
  //: IN g2 (D) @(192,114) /sn:0 /w:[ 5 ]
  INV1 g1 (.in(D), .out(w0));   //: @(269, 124) /sz:(40, 40) /sn:0 /p:[ Li0>0 Ro0<1 ]
  //: OUT g5 (Y) @(424,125) /sn:0 /w:[ 1 ]
  FFSR g0 (.S(D), .R(w0), .clk(Clk), .Y(Y));   //: @(357, 107) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>0 Bi0>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin REG4
module REG4(out, Clk, in);
//: interface  /sz:(75, 52) /bd:[ Ti0>Clk(37/75) Li0>in[3:0](25/52) Ro0<out[3:0](25/52) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] in;    //: /sn:0 {0}(#:148,-71)(148,-19){1}
//: {2}(148,-18)(148,55){3}
//: {4}(148,56)(148,130){5}
//: {6}(148,131)(148,202){7}
//: {8}(148,203)(148,213){9}
input Clk;    //: /sn:0 {0}(202,-73)(202,14){1}
//: {2}(204,16)(261,16)(261,4){3}
//: {4}(202,18)(202,83){5}
//: {6}(204,85)(259,85)(259,78){7}
//: {8}(202,87)(202,157){9}
//: {10}(204,159)(260,159)(260,153){11}
//: {12}(202,161)(202,236)(260,236)(260,225){13}
output [3:0] out;    //: /sn:0 {0}(#:454,212)(494,212){1}
wire w6;    //: /sn:0 {0}(152,131)(241,131){1}
wire w3;    //: /sn:0 {0}(152,56)(240,56){1}
wire w0;    //: /sn:0 {0}(152,-18)(242,-18){1}
wire w8;    //: /sn:0 {0}(283,131)(399,131)(399,217)(448,217){1}
wire w2;    //: /sn:0 {0}(284,-18)(418,-18)(418,197)(448,197){1}
wire w11;    //: /sn:0 {0}(283,203)(309,203)(309,227)(448,227){1}
wire w5;    //: /sn:0 {0}(282,56)(409,56)(409,207)(448,207){1}
wire w9;    //: /sn:0 {0}(152,203)(241,203){1}
//: enddecls

  FFD g4 (.D(w3), .Clk(Clk), .Y(w5));   //: @(241, 37) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>7 Ro0<0 ]
  //: joint g8 (Clk) @(202, 159) /w:[ 10 9 -1 12 ]
  FFD g3 (.D(w0), .Clk(Clk), .Y(w2));   //: @(243, -37) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>3 Ro0<0 ]
  assign w0 = in[0]; //: TAP g17 @(146,-18) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: OUT g2 (out) @(491,212) /sn:0 /w:[ 1 ]
  assign out = {w11, w8, w5, w2}; //: CONCAT g1  @(453,212) /sn:0 /w:[ 0 1 1 1 1 ] /dr:1 /tp:1 /drp:1
  assign w3 = in[1]; //: TAP g18 @(146,56) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g10 (Clk) @(202, 16) /w:[ 2 1 -1 4 ]
  FFD g6 (.D(w9), .Clk(Clk), .Y(w11));   //: @(242, 184) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>13 Ro0<0 ]
  //: IN g7 (Clk) @(202,-75) /sn:0 /R:3 /w:[ 0 ]
  //: joint g9 (Clk) @(202, 85) /w:[ 6 5 -1 8 ]
  FFD g5 (.D(w6), .Clk(Clk), .Y(w8));   //: @(242, 112) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>11 Ro0<0 ]
  assign w6 = in[2]; //: TAP g19 @(146,131) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  assign w9 = in[3]; //: TAP g20 @(146,203) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: IN g0 (in) @(148,-73) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin AND2
module AND2(in2, in1, out);
//: interface  /sz:(40, 40) /bd:[ Li0>in2(30/40) Li1>in1(10/40) Ro0<out(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input in1;    //: /sn:0 {0}(275,165)(201,165)(201,154)(186,154){1}
output out;    //: /sn:0 {0}(410,175)(443,175){1}
input in2;    //: /sn:0 {0}(275,185)(199,185)(199,193)(184,193){1}
wire w0;    //: /sn:0 {0}(317,173)(368,173){1}
//: enddecls

  //: IN g4 (in2) @(182,193) /sn:0 /w:[ 1 ]
  //: IN g3 (in1) @(184,154) /sn:0 /w:[ 1 ]
  //: OUT g2 (out) @(440,175) /sn:0 /w:[ 1 ]
  INV1 g1 (.in(w0), .out(out));   //: @(369, 155) /sz:(40, 40) /sn:0 /p:[ Li0>1 Ro0<0 ]
  NAND2 g0 (.in1(in1), .in2(in2), .out(w0));   //: @(276, 155) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX2
module MUX2(out, c, in0, in1);
//: interface  /sz:(68, 72) /bd:[ Li0>in0(16/72) Li1>in1(48/72) Bi0>c(30/68) Ro0<out(32/72) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input in1;    //: /sn:0 {0}(75,207)(221,207){1}
input in0;    //: /sn:0 {0}(78,88)(225,88){1}
output out;    //: /sn:0 {0}(381,155)(410,155){1}
input c;    //: /sn:0 {0}(153,275)(153,229){1}
//: {2}(155,227)(221,227){3}
//: {4}(153,225)(153,183){5}
wire w1;    //: /sn:0 {0}(152,141)(152,108)(225,108){1}
wire w2;    //: /sn:0 {0}(267,96)(324,96)(324,147)(339,147){1}
wire w5;    //: /sn:0 {0}(263,215)(324,215)(324,167)(339,167){1}
//: enddecls

  //: OUT g8 (out) @(407,155) /sn:0 /w:[ 1 ]
  //: IN g4 (c) @(153,277) /sn:0 /R:1 /w:[ 0 ]
  INV1 g3 (.in(c), .out(w1));   //: @(132, 142) /sz:(40, 40) /R:1 /sn:0 /p:[ Bi0>5 To0<0 ]
  NAND2 g2 (.in2(w5), .in1(w2), .out(out));   //: @(340, 137) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  NAND2 g1 (.in2(c), .in1(in1), .out(w5));   //: @(222, 197) /sz:(40, 40) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]
  //: IN g6 (in0) @(76,88) /sn:0 /w:[ 0 ]
  //: IN g7 (in1) @(73,207) /sn:0 /w:[ 0 ]
  //: joint g5 (c) @(153, 227) /w:[ 2 4 -1 1 ]
  NAND2 g0 (.in2(w1), .in1(in0), .out(w2));   //: @(226, 78) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FFD
module FFD(Clk, Y, D);
//: interface  /sz:(40, 40) /bd:[ Li0>D(19/40) Bi0>Clk(18/40) Ro0<Y(19/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(375,157)(416,157){1}
//: {2}(418,155)(418,124){3}
//: {4}(418,159)(418,189){5}
input D;    //: /sn:0 {0}(238,102)(278,102){1}
output Y;    //: /sn:0 {0}(441,102)(485,102){1}
wire w1;    //: /sn:0 {0}(333,158)(297,158)(297,124){1}
wire w2;    //: /sn:0 {0}(320,102)(399,102){1}
//: enddecls

  //: joint g4 (Clk) @(418, 157) /w:[ -1 2 1 4 ]
  INV1 g3 (.in(Clk), .out(w1));   //: @(334, 138) /sz:(40, 40) /R:2 /sn:0 /p:[ Ri0>0 Lo0<0 ]
  //: IN g2 (Clk) @(418,191) /sn:0 /R:1 /w:[ 5 ]
  FFDLS g1 (.D(w2), .Clk(Clk), .Y(Y));   //: @(400, 83) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>3 Ro0<0 ]
  //: OUT g6 (Y) @(482,102) /sn:0 /w:[ 1 ]
  //: IN g5 (D) @(236,102) /sn:0 /w:[ 0 ]
  FFDLS g0 (.D(D), .Clk(w1), .Y(w2));   //: @(279, 83) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin INV1
module INV1(in, out);
//: interface  /sz:(40, 40) /bd:[ Li0>in(21/40) Ro0<out(20/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply1 w6;    //: /sn:0 {0}(320,95)(320,123){1}
input in;    //: /sn:0 {0}(254,164)(289,164){1}
//: {2}(291,162)(291,131)(306,131){3}
//: {4}(291,166)(291,200)(306,200){5}
supply0 w3;    //: /sn:0 {0}(320,209)(320,234){1}
output out;    //: /sn:0 {0}(320,140)(320,161){1}
//: {2}(322,163)(359,163){3}
//: {4}(320,165)(320,192){5}
//: enddecls

  //: IN g4 (in) @(252,164) /sn:0 /w:[ 0 ]
  //: VDD g3 (w6) @(331,95) /sn:0 /w:[ 0 ]
  //: GROUND g2 (w3) @(320,240) /sn:0 /w:[ 1 ]
  _GGNMOS #(2, 1) g1 (.Z(out), .S(w3), .G(in));   //: @(314,200) /sn:0 /w:[ 5 0 5 ]
  //: joint g6 (in) @(291, 164) /w:[ -1 2 1 4 ]
  //: joint g7 (out) @(320, 163) /w:[ 2 1 -1 4 ]
  //: OUT g5 (out) @(356,163) /sn:0 /w:[ 3 ]
  _GGPMOS #(2, 1) g0 (.Z(out), .S(w6), .G(in));   //: @(314,131) /sn:0 /w:[ 0 1 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin NAND2
module NAND2(in1, out, in2);
//: interface  /sz:(40, 40) /bd:[ Li0>in1(10/40) Li1>in2(30/40) Ro0<out(18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w6;    //: /sn:0 {0}(154,1)(154,18){1}
//: {2}(156,20)(184,20)(184,26){3}
//: {4}(152,20)(127,20)(127,42){5}
supply0 w3;    //: /sn:0 {0}(155,184)(155,222){1}
input in1;    //: /sn:0 {0}(47,34)(73,34){1}
//: {2}(77,34)(170,34){3}
//: {4}(75,36)(75,117)(141,117){5}
output out;    //: /sn:0 {0}(155,109)(155,90){1}
//: {2}(157,88)(214,88){3}
//: {4}(155,86)(155,76){5}
//: {6}(157,74)(184,74)(184,43){7}
//: {8}(153,74)(127,74)(127,59){9}
input in2;    //: /sn:0 {0}(52,126)(101,126){1}
//: {2}(103,124)(103,50)(113,50){3}
//: {4}(103,128)(103,175)(141,175){5}
wire w4;    //: /sn:0 {0}(155,126)(155,167){1}
//: enddecls

  //: IN g8 (in1) @(45,34) /sn:0 /w:[ 0 ]
  //: joint g4 (out) @(155, 74) /w:[ 6 -1 8 5 ]
  _GGNMOS #(2, 1) g3 (.Z(w4), .S(w3), .G(in2));   //: @(149,175) /sn:0 /w:[ 1 0 5 ]
  _GGPMOS #(2, 1) g2 (.Z(out), .S(w6), .G(in1));   //: @(178,34) /sn:0 /w:[ 7 3 3 ]
  _GGNMOS #(2, 1) g1 (.Z(out), .S(w4), .G(in1));   //: @(149,117) /sn:0 /w:[ 0 0 5 ]
  //: OUT g10 (out) @(211,88) /sn:0 /w:[ 3 ]
  //: VDD g6 (w6) @(165,1) /sn:0 /w:[ 0 ]
  //: IN g9 (in2) @(50,126) /sn:0 /w:[ 0 ]
  //: joint g7 (w6) @(154, 20) /w:[ 2 1 4 -1 ]
  //: joint g12 (in1) @(75, 34) /w:[ 2 -1 1 4 ]
  //: joint g11 (out) @(155, 88) /w:[ 2 4 -1 1 ]
  //: GROUND g5 (w3) @(155,228) /sn:0 /w:[ 1 ]
  _GGPMOS #(2, 1) g0 (.Z(out), .S(w6), .G(in2));   //: @(121,50) /sn:0 /w:[ 9 5 3 ]
  //: joint g13 (in2) @(103, 126) /w:[ -1 2 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin MUX8
module MUX8(a, C, b, out);
//: interface  /sz:(40, 50) /bd:[ Ti0>C(19/40) Li0>a[7:0](12/50) Li1>b[7:0](38/50) Ro0<out[7:0](24/50) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] b;    //: /sn:0 {0}(#:7,45)(79,45){1}
//: {2}(80,45)(198,45){3}
//: {4}(199,45)(313,45){5}
//: {6}(314,45)(437,45){7}
//: {8}(438,45)(556,45){9}
//: {10}(557,45)(671,45){11}
//: {12}(672,45)(799,45){13}
//: {14}(800,45)(914,45){15}
//: {16}(915,45)(#:921,45){17}
output [7:0] out;    //: /sn:0 {0}(#:512,343)(512,379){1}
input C;    //: /sn:0 {0}(174,171)(158,171)(158,98){1}
//: {2}(160,96)(271,96){3}
//: {4}(275,96)(393,96){5}
//: {6}(397,96)(515,96){7}
//: {8}(519,96)(625,96){9}
//: {10}(629,96)(761,96){11}
//: {12}(765,96)(869,96){13}
//: {14}(873,96)(975,96){15}
//: {16}(871,98)(871,178)(890,178){17}
//: {18}(763,98)(763,176)(775,176){19}
//: {20}(627,98)(627,176)(647,176){21}
//: {22}(517,98)(517,174)(532,174){23}
//: {24}(395,98)(395,175)(413,175){25}
//: {26}(273,98)(273,173)(289,173){27}
//: {28}(156,96)(40,96)(40,172)(55,172){29}
input [7:0] a;    //: /sn:0 {0}(#:8,15)(111,15){1}
//: {2}(112,15)(230,15){3}
//: {4}(231,15)(345,15){5}
//: {6}(346,15)(469,15){7}
//: {8}(470,15)(588,15){9}
//: {10}(589,15)(703,15){11}
//: {12}(704,15)(831,15){13}
//: {14}(832,15)(946,15){15}
//: {16}(947,15)(954,15){17}
wire w6;    //: /sn:0 {0}(487,337)(487,305)(215,305)(215,210){1}
wire w16;    //: /sn:0 {0}(557,143)(557,49){1}
wire w13;    //: /sn:0 {0}(704,145)(704,19){1}
wire w25;    //: /sn:0 {0}(947,147)(947,19){1}
wire w4;    //: /sn:0 {0}(231,140)(231,19){1}
wire w22;    //: /sn:0 {0}(527,337)(527,295)(688,295)(688,215){1}
wire w3;    //: /sn:0 {0}(477,337)(477,315)(96,315)(96,211){1}
wire w0;    //: /sn:0 {0}(112,141)(112,19){1}
wire w20;    //: /sn:0 {0}(438,144)(438,49){1}
wire w30;    //: /sn:0 {0}(547,337)(547,313)(931,313)(931,217){1}
wire w29;    //: /sn:0 {0}(832,145)(832,19){1}
wire w18;    //: /sn:0 {0}(517,337)(517,287)(573,287)(573,213){1}
wire w12;    //: /sn:0 {0}(672,145)(672,49){1}
wire w10;    //: /sn:0 {0}(497,337)(497,296)(330,296)(330,212){1}
wire w23;    //: /sn:0 {0}(507,337)(507,288)(454,288)(454,214){1}
wire w24;    //: /sn:0 {0}(314,142)(314,49){1}
wire w21;    //: /sn:0 {0}(470,144)(470,19){1}
wire w31;    //: /sn:0 {0}(816,215)(816,302)(537,302)(537,337){1}
wire w1;    //: /sn:0 {0}(80,141)(80,49){1}
wire w32;    //: /sn:0 {0}(915,147)(915,49){1}
wire w8;    //: /sn:0 {0}(346,142)(346,19){1}
wire w17;    //: /sn:0 {0}(589,143)(589,19){1}
wire w28;    //: /sn:0 {0}(800,145)(800,49){1}
wire w5;    //: /sn:0 {0}(199,140)(199,49){1}
//: enddecls

  MUX2 g8 (.in1(w28), .in0(w29), .c(C), .out(w31));   //: @(776, 146) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>19 Bo0<0 ]
  MUX2 g4 (.in1(w12), .in0(w13), .c(C), .out(w22));   //: @(648, 146) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>21 Bo0<1 ]
  assign w28 = b[1]; //: TAP g16 @(800,43) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  //: IN g3 (a) @(6,15) /sn:0 /w:[ 0 ]
  //: IN g26 (C) @(977,96) /sn:0 /R:2 /w:[ 15 ]
  assign w32 = b[0]; //: TAP g17 @(915,43) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  MUX2 g2 (.in1(w24), .in0(w8), .c(C), .out(w10));   //: @(290, 143) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>27 Bo0<1 ]
  //: joint g30 (C) @(517, 96) /w:[ 8 -1 7 22 ]
  assign w13 = a[2]; //: TAP g23 @(704,13) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  assign w29 = a[1]; //: TAP g24 @(832,13) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  MUX2 g1 (.in1(w5), .in0(w4), .c(C), .out(w6));   //: @(175, 141) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 ]
  //: joint g29 (C) @(627, 96) /w:[ 10 -1 9 20 ]
  assign w0 = a[7]; //: TAP g18 @(112,13) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w25 = a[0]; //: TAP g25 @(947,13) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  assign w1 = b[7]; //: TAP g10 @(80,43) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  MUX2 g6 (.in1(w20), .in0(w21), .c(C), .out(w23));   //: @(414, 145) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>25 Bo0<1 ]
  //: IN g9 (b) @(5,45) /sn:0 /w:[ 0 ]
  MUX2 g7 (.in1(w32), .in0(w25), .c(C), .out(w30));   //: @(891, 148) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>17 Bo0<1 ]
  //: OUT g35 (out) @(512,376) /sn:0 /R:3 /w:[ 1 ]
  //: joint g31 (C) @(395, 96) /w:[ 6 -1 5 24 ]
  assign w17 = a[3]; //: TAP g22 @(589,13) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  //: joint g33 (C) @(158, 96) /w:[ 2 -1 28 1 ]
  assign w24 = b[5]; //: TAP g12 @(314,43) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign out = {w3, w6, w10, w23, w18, w22, w31, w30}; //: CONCAT g34  @(512,342) /sn:0 /R:3 /w:[ 0 0 0 0 0 0 0 1 0 ] /dr:0 /tp:0 /drp:1
  //: joint g28 (C) @(763, 96) /w:[ 12 -1 11 18 ]
  assign w16 = b[3]; //: TAP g14 @(557,43) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign w5 = b[6]; //: TAP g11 @(199,43) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  MUX2 g5 (.in1(w16), .in0(w17), .c(C), .out(w18));   //: @(533, 144) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>23 Bo0<1 ]
  assign w21 = a[4]; //: TAP g21 @(470,13) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w4 = a[6]; //: TAP g19 @(231,13) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: joint g32 (C) @(273, 96) /w:[ 4 -1 3 26 ]
  assign w8 = a[5]; //: TAP g20 @(346,13) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign w12 = b[2]; //: TAP g15 @(672,43) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  MUX2 g0 (.in1(w1), .in0(w0), .c(C), .out(w3));   //: @(56, 142) /sz:(72, 68) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Li0>29 Bo0<1 ]
  //: joint g27 (C) @(871, 96) /w:[ 14 -1 13 16 ]
  assign w20 = b[4]; //: TAP g13 @(438,43) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin NOR2
module NOR2(in1, out, in2);
//: interface  /sz:(40, 40) /bd:[ Li0>in2(30/40) Li1>in1(8/40) Ro0<out(18/40) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w0;    //: /sn:0 {0}(270,113)(270,137){1}
input in1;    //: /sn:0 {0}(129,145)(189,145){1}
//: {2}(193,145)(256,145){3}
//: {4}(191,147)(191,287)(292,287){5}
supply0 w1;    //: /sn:0 {0}(269,356)(269,332){1}
//: {2}(271,330)(306,330)(306,296){3}
//: {4}(267,330)(235,330)(235,319){5}
output out;    //: /sn:0 {0}(270,219)(270,235){1}
//: {2}(272,237)(371,237){3}
//: {4}(270,239)(270,270){5}
//: {6}(272,272)(306,272)(306,279){7}
//: {8}(268,272)(235,272)(235,302){9}
input in2;    //: /sn:0 {0}(126,210)(157,210){1}
//: {2}(161,210)(256,210){3}
//: {4}(159,212)(159,310)(221,310){5}
wire w2;    //: /sn:0 {0}(270,154)(270,202){1}
//: enddecls

  _GGNMOS #(2, 1) g4 (.Z(out), .S(w1), .G(in2));   //: @(229,310) /sn:0 /w:[ 9 5 5 ]
  //: IN g8 (in1) @(127,145) /sn:0 /w:[ 0 ]
  _GGPMOS #(2, 1) g3 (.Z(out), .S(w2), .G(in2));   //: @(264,210) /sn:0 /w:[ 0 1 3 ]
  _GGPMOS #(2, 1) g2 (.Z(w2), .S(w0), .G(in1));   //: @(264,145) /sn:0 /w:[ 0 1 3 ]
  //: GROUND g1 (w1) @(269,362) /sn:0 /w:[ 0 ]
  //: OUT g10 (out) @(368,237) /sn:0 /w:[ 3 ]
  //: joint g6 (w1) @(269, 330) /w:[ 2 -1 4 1 ]
  //: joint g7 (out) @(270, 272) /w:[ 6 5 8 -1 ]
  //: IN g9 (in2) @(124,210) /sn:0 /w:[ 0 ]
  //: joint g12 (in1) @(191, 145) /w:[ 2 -1 1 4 ]
  //: joint g11 (out) @(270, 237) /w:[ 2 1 -1 4 ]
  _GGNMOS #(2, 1) g5 (.Z(out), .S(w1), .G(in1));   //: @(300,287) /sn:0 /w:[ 7 3 5 ]
  //: VDD g0 (w0) @(281,113) /sn:0 /w:[ 0 ]
  //: joint g13 (in2) @(159, 210) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA12
module FA12(cin, s, cout, b, a);
//: interface  /sz:(77, 74) /bd:[ Ti0>b[11:0](54/77) Ti1>a[11:0](15/77) Ri0>cin(36/74) Lo0<cout(34/74) Bo0<s[11:0](35/77) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [11:0] b;    //: /sn:0 {0}(#:402,168)(405,168){1}
//: {2}(406,168)(420,168){3}
//: {4}(421,168)(434,168){5}
//: {6}(435,168)(450,168){7}
//: {8}(451,168)(965,168){9}
//: {10}(966,168)(985,168){11}
//: {12}(986,168)(1004,168){13}
//: {14}(1005,168)(1022,168){15}
//: {16}(1023,168)(1040,168){17}
//: {18}(1041,168)(1059,168){19}
//: {20}(1060,168)(1075,168){21}
//: {22}(1076,168)(1093,168){23}
//: {24}(1094,168)(#:1214,168){25}
input cin;    //: /sn:0 {0}(1225,387)(955,387){1}
output [11:0] s;    //: /sn:0 {0}(#:660,504)(660,541){1}
output cout;    //: /sn:0 {0}(339,380)(279,380){1}
input [11:0] a;    //: /sn:0 {0}(#:286,76)(289,76){1}
//: {2}(290,76)(304,76){3}
//: {4}(305,76)(318,76){5}
//: {6}(319,76)(334,76){7}
//: {8}(335,76)(670,76){9}
//: {10}(671,76)(688,76){11}
//: {12}(689,76)(706,76){13}
//: {14}(707,76)(722,76){15}
//: {16}(723,76)(739,76){17}
//: {18}(740,76)(754,76){19}
//: {20}(755,76)(769,76){21}
//: {22}(770,76)(786,76){23}
//: {24}(787,76)(#:1206,76){25}
wire w16;    //: /sn:0 {0}(966,172)(966,249)(1024,249)(1024,283){1}
wire w13;    //: /sn:0 {0}(1054,283)(1054,217)(1023,217)(1023,172){1}
wire w6;    //: /sn:0 {0}(1084,283)(1084,193)(1076,193)(1076,172){1}
wire w7;    //: /sn:0 {0}(1074,283)(1074,200)(1060,200)(1060,172){1}
wire [3:0] w34;    //: /sn:0 {0}(#:320,294)(320,344)(359,344)(#:359,359){1}
wire w4;    //: /sn:0 {0}(757,291)(757,118)(740,118)(740,80){1}
wire [7:0] w22;    //: /sn:0 {0}(665,498)(665,432)(#:917,432)(#:917,422){1}
wire w3;    //: /sn:0 {0}(767,291)(767,110)(755,110)(755,80){1}
wire w0;    //: /sn:0 {0}(1094,172)(1094,283){1}
wire w20;    //: /sn:0 {0}(420,388)(884,388){1}
wire [3:0] w29;    //: /sn:0 {0}(655,498)(655,432)(#:385,432)(#:385,412){1}
wire w30;    //: /sn:0 {0}(315,288)(315,106)(305,106)(305,80){1}
wire [3:0] w18;    //: /sn:0 {0}(#:436,296)(436,344)(395,344)(#:395,359){1}
wire w19;    //: /sn:0 {0}(737,291)(737,139)(707,139)(707,80){1}
wire w12;    //: /sn:0 {0}(717,291)(717,160)(671,160)(671,80){1}
wire w23;    //: /sn:0 {0}(431,290)(431,198)(421,198)(421,172){1}
wire w10;    //: /sn:0 {0}(435,172)(435,188)(441,188)(441,290){1}
wire w24;    //: /sn:0 {0}(421,290)(421,209)(406,209)(406,172){1}
wire w21;    //: /sn:0 {0}(747,291)(747,127)(723,127)(723,80){1}
wire w31;    //: /sn:0 {0}(335,80)(335,288){1}
wire w1;    //: /sn:0 {0}(770,80)(770,102)(777,102)(777,291){1}
wire w32;    //: /sn:0 {0}(319,80)(319,96)(325,96)(325,288){1}
wire w8;    //: /sn:0 {0}(1064,283)(1064,208)(1041,208)(1041,172){1}
wire [7:0] w17;    //: /sn:0 {0}(#:752,297)(752,340)(#:899,340)(#:899,355){1}
wire w33;    //: /sn:0 {0}(305,288)(305,117)(290,117)(290,80){1}
wire w14;    //: /sn:0 {0}(1044,283)(1044,228)(1005,228)(1005,172){1}
wire w11;    //: /sn:0 {0}(727,291)(727,150)(689,150)(689,80){1}
wire [7:0] w2;    //: /sn:0 {0}(#:1059,289)(1059,340)(#:932,340)(#:932,355){1}
wire w15;    //: /sn:0 {0}(986,172)(986,238)(1034,238)(1034,283){1}
wire w5;    //: /sn:0 {0}(451,172)(451,290){1}
wire w9;    //: /sn:0 {0}(787,80)(787,291){1}
//: enddecls

  assign w6 = b[1]; //: TAP g8 @(1076,166) /sn:0 /R:1 /w:[ 1 21 22 ] /ss:1
  assign w1 = a[1]; //: TAP g4 @(770,74) /sn:0 /R:1 /w:[ 0 21 22 ] /ss:1
  assign w21 = a[4]; //: TAP g16 @(723,74) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  assign w9 = a[0]; //: TAP g3 @(787,74) /sn:0 /R:1 /w:[ 0 23 24 ] /ss:1
  assign w23 = b[10]; //: TAP g26 @(421,166) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w19 = a[5]; //: TAP g17 @(707,74) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  assign w2 = {w16, w15, w14, w13, w8, w7, w6, w0}; //: CONCAT g2  @(1059,288) /sn:0 /R:3 /w:[ 0 1 1 0 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  FA4 g23 (.a(w34), .b(w18), .cin(w20), .cout(cout), .s(w29));   //: @(340, 360) /sz:(79, 51) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<1 ]
  assign w32 = a[9]; //: TAP g30 @(319,74) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w5 = b[8]; //: TAP g24 @(451,166) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: IN g1 (cin) @(1227,387) /sn:0 /R:2 /w:[ 0 ]
  assign w31 = a[8]; //: TAP g29 @(335,74) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w11 = a[6]; //: TAP g18 @(689,74) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  assign w10 = b[9]; //: TAP g25 @(435,166) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w8 = b[3]; //: TAP g10 @(1041,166) /sn:0 /R:1 /w:[ 1 17 18 ] /ss:1
  assign w4 = a[3]; //: TAP g6 @(740,74) /sn:0 /R:1 /w:[ 1 17 18 ] /ss:1
  //: OUT g35 (s) @(660,538) /sn:0 /R:3 /w:[ 1 ]
  assign w7 = b[2]; //: TAP g9 @(1060,166) /sn:0 /R:1 /w:[ 1 19 20 ] /ss:1
  assign w0 = b[0]; //: TAP g7 @(1094,166) /sn:0 /R:1 /w:[ 0 23 24 ] /ss:1
  assign w34 = {w33, w30, w32, w31}; //: CONCAT g31  @(320,293) /sn:0 /R:3 /w:[ 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  assign w18 = {w24, w23, w10, w5}; //: CONCAT g22  @(436,295) /sn:0 /R:3 /w:[ 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g33 (cout) @(282,380) /sn:0 /R:2 /w:[ 1 ]
  assign w13 = b[4]; //: TAP g12 @(1023,166) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  assign s = {w29, w22}; //: CONCAT g34  @(660,503) /sn:0 /R:3 /w:[ 0 0 0 ] /dr:1 /tp:0 /drp:1
  assign w30 = a[10]; //: TAP g28 @(305,74) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w15 = b[6]; //: TAP g14 @(986,166) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  assign w3 = a[2]; //: TAP g11 @(755,74) /sn:0 /R:1 /w:[ 1 19 20 ] /ss:1
  //: IN g5 (b) @(1216,168) /sn:0 /R:2 /w:[ 25 ]
  assign w14 = b[5]; //: TAP g21 @(1005,166) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  assign w12 = a[7]; //: TAP g19 @(671,74) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign w33 = a[11]; //: TAP g32 @(290,74) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w16 = b[7]; //: TAP g20 @(966,166) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  FA8 g0 (.a(w17), .b(w2), .cin(cin), .cout(w20), .s(w22));   //: @(885, 356) /sz:(69, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  //: IN g15 (a) @(1208,76) /sn:0 /R:2 /w:[ 25 ]
  assign w24 = b[11]; //: TAP g27 @(406,166) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w17 = {w12, w11, w19, w21, w4, w3, w1, w9}; //: CONCAT g13  @(752,296) /sn:0 /R:3 /w:[ 0 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1

endmodule
//: /netlistEnd

//: /netlistBegin MUL8
module MUL8(b, out, a);
//: interface  /sz:(63, 62) /bd:[ Li0>a[7:0](14/62) Li1>b[7:0](44/62) Ro0<out[15:0](32/62) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
supply0 [2:0] w58;    //: /sn:0 {0}(#:709,706)(#:709,785){1}
input [7:0] b;    //: /sn:0 {0}(#:101,173)(106,173){1}
//: {2}(107,173)(124,173){3}
//: {4}(125,173)(144,173){5}
//: {6}(145,173)(160,173){7}
//: {8}(161,173)(414,173){9}
//: {10}(415,173)(432,173){11}
//: {12}(433,173)(451,173){13}
//: {14}(452,173)(467,173){15}
//: {16}(468,173)(705,173){17}
//: {18}(706,173)(723,173){19}
//: {20}(724,173)(743,173){21}
//: {22}(744,173)(759,173){23}
//: {24}(760,173)(1013,173){25}
//: {26}(1014,173)(1031,173){27}
//: {28}(1032,173)(1050,173){29}
//: {30}(1051,173)(1066,173){31}
//: {32}(1067,173)(#:1227,173){33}
supply0 w72;    //: /sn:0 {0}(690,871)(656,871){1}
supply0 w56;    //: /sn:0 {0}(956,693)(928,693){1}
supply0 w71;    //: /sn:0 {0}(260,705)(224,705){1}
supply0 w70;    //: /sn:0 {0}(359,704)(331,704){1}
output [15:0] out;    //: /sn:0 {0}(#:1095,996)(1095,1038){1}
supply0 [3:0] w67;    //: /sn:0 {0}(#:427,555)(#:427,632){1}
input [7:0] a;    //: /sn:0 {0}(#:148,81)(152,81){1}
//: {2}(153,81)(169,81){3}
//: {4}(170,81)(184,81){5}
//: {6}(185,81)(200,81){7}
//: {8}(201,81)(459,81){9}
//: {10}(460,81)(477,81){11}
//: {12}(478,81)(493,81){13}
//: {14}(494,81)(507,81){15}
//: {16}(508,81)(751,81){17}
//: {18}(752,81)(768,81){19}
//: {20}(769,81)(783,81){21}
//: {22}(784,81)(799,81){23}
//: {24}(800,81)(1058,81){25}
//: {26}(1059,81)(1076,81){27}
//: {28}(1077,81)(1092,81){29}
//: {30}(1093,81)(1106,81){31}
//: {32}(1107,81)(#:1219,81){33}
supply0 w77;    //: /sn:0 {0}(541,869)(577,869){1}
supply0 [3:0] w40;    //: /sn:0 {0}(#:1026,545)(#:1026,622){1}
wire w16;    //: /sn:0 {0}(730,296)(730,220)(706,220)(706,177){1}
wire w13;    //: /sn:0 {0}(760,296)(760,177){1}
wire w6;    //: /sn:0 {0}(1057,288)(1057,197)(1051,197)(1051,177){1}
wire w65;    //: /sn:0 {0}(447,521)(447,632){1}
wire w7;    //: /sn:0 {0}(1047,288)(1047,208)(1032,208)(1032,177){1}
wire w50;    //: /sn:0 {0}(1076,511)(1076,606)(1085,606)(1085,990){1}
wire w34;    //: /sn:0 {0}(131,296)(131,220)(107,220)(107,177){1}
wire w59;    //: /sn:0 {0}(467,521)(467,632){1}
wire [11:0] w62;    //: /sn:0 {0}(632,834)(632,806)(#:719,806)(#:719,791){1}
wire [3:0] w39;    //: /sn:0 {0}(770,344)(770,379)(#:777,379)(777,394){1}
wire w25;    //: /sn:0 {0}(468,288)(468,177){1}
wire w4;    //: /sn:0 {0}(1077,288)(1077,132)(1059,132)(1059,85){1}
wire [3:0] w36;    //: /sn:0 {0}(1077,343)(1077,378)(#:1084,378)(1084,393){1}
wire w22;    //: /sn:0 {0}(185,85)(185,110)(191,110)(191,296){1}
wire w3;    //: /sn:0 {0}(1087,288)(1087,118)(1077,118)(1077,85){1}
wire w0;    //: /sn:0 {0}(1107,85)(1107,288){1}
wire w60;    //: /sn:0 {0}(857,694)(719,694)(719,785){1}
wire w20;    //: /sn:0 {0}(508,85)(508,288){1}
wire w30;    //: /sn:0 {0}(161,296)(161,177){1}
wire w29;    //: /sn:0 {0}(181,296)(181,116)(170,116)(170,85){1}
wire [3:0] w42;    //: /sn:0 {0}(468,336)(468,371)(#:461,371)(461,386){1}
wire [3:0] w37;    //: /sn:0 {0}(1067,343)(1067,378)(#:1060,378)(1060,393){1}
wire w73;    //: /sn:0 {0}(507,521)(507,589)(519,589)(519,786){1}
wire w66;    //: /sn:0 {0}(437,521)(437,632){1}
wire w19;    //: /sn:0 {0}(458,288)(458,197)(452,197)(452,177){1}
wire w18;    //: /sn:0 {0}(494,85)(494,115)(498,115)(498,288){1}
wire w12;    //: /sn:0 {0}(770,296)(770,130)(752,130)(752,85){1}
wire w63;    //: /sn:0 {0}(457,521)(457,632){1}
wire w23;    //: /sn:0 {0}(488,288)(488,118)(478,118)(478,85){1}
wire w10;    //: /sn:0 {0}(784,85)(784,110)(790,110)(790,296){1}
wire [7:0] w54;    //: /sn:0 {0}(#:1071,505)(1071,451){1}
wire w24;    //: /sn:0 {0}(478,288)(478,132)(460,132)(460,85){1}
wire w21;    //: /sn:0 {0}(201,85)(201,296){1}
wire w31;    //: /sn:0 {0}(171,296)(171,130)(153,130)(153,85){1}
wire w1;    //: /sn:0 {0}(1093,85)(1093,115)(1097,115)(1097,288){1}
wire [7:0] w68;    //: /sn:0 {0}(#:447,638)(447,651)(#:308,651)(#:308,672){1}
wire w32;    //: /sn:0 {0}(151,296)(151,195)(145,195)(145,177){1}
wire w53;    //: /sn:0 {0}(1046,511)(1046,622){1}
wire [3:0] w46;    //: /sn:0 {0}(171,337)(171,372)(#:178,372)(178,387){1}
wire w8;    //: /sn:0 {0}(1037,288)(1037,222)(1014,222)(1014,177){1}
wire w52;    //: /sn:0 {0}(1056,511)(1056,622){1}
wire w75;    //: /sn:0 {0}(487,521)(487,611)(499,611)(499,786){1}
wire [7:0] w44;    //: /sn:0 {0}(#:472,515)(472,444){1}
wire w27;    //: /sn:0 {0}(438,288)(438,222)(415,222)(415,177){1}
wire [7:0] w17;    //: /sn:0 {0}(#:765,338)(#:765,302){1}
wire [7:0] w35;    //: /sn:0 {0}(#:166,331)(#:166,302){1}
wire w33;    //: /sn:0 {0}(141,296)(141,206)(125,206)(125,177){1}
wire [7:0] w28;    //: /sn:0 {0}(#:473,330)(#:473,294){1}
wire [7:0] w69;    //: /sn:0 {0}(#:293,739)(293,771)(#:479,771)(#:479,786){1}
wire w49;    //: /sn:0 {0}(1096,511)(1096,591)(1105,591)(1105,990){1}
wire [3:0] w45;    //: /sn:0 {0}(161,337)(161,372)(#:154,372)(154,387){1}
wire w14;    //: /sn:0 {0}(750,296)(750,195)(744,195)(744,177){1}
wire [11:0] w78;    //: /sn:0 {0}(593,834)(593,807)(#:499,807)(#:499,792){1}
wire w74;    //: /sn:0 {0}(497,521)(497,602)(509,602)(509,786){1}
wire w48;    //: /sn:0 {0}(1106,511)(1106,580)(1115,580)(1115,990){1}
wire [7:0] w41;    //: /sn:0 {0}(764,452)(764,646)(#:872,646)(#:872,661){1}
wire w11;    //: /sn:0 {0}(780,296)(780,116)(769,116)(769,85){1}
wire [7:0] w2;    //: /sn:0 {0}(#:1072,294)(#:1072,337){1}
wire [7:0] w47;    //: /sn:0 {0}(#:275,672)(#:275,654)(165,654)(165,445){1}
wire [11:0] w83;    //: /sn:0 {0}(613,910)(613,943)(1075,943)(#:1075,990){1}
wire w15;    //: /sn:0 {0}(740,296)(740,206)(724,206)(724,177){1}
wire [7:0] w61;    //: /sn:0 {0}(729,785)(729,743)(#:890,743)(#:890,728){1}
wire w55;    //: /sn:0 {0}(1086,511)(1086,600)(1095,600)(1095,990){1}
wire [3:0] w38;    //: /sn:0 {0}(760,344)(760,379)(#:753,379)(753,394){1}
wire w5;    //: /sn:0 {0}(1067,288)(1067,177){1}
wire [7:0] w64;    //: /sn:0 {0}(#:1046,628)(1046,641)(#:905,641)(#:905,661){1}
wire [3:0] w43;    //: /sn:0 {0}(478,336)(478,371)(#:485,371)(485,386){1}
wire w76;    //: /sn:0 {0}(477,521)(477,622)(489,622)(489,786){1}
wire w26;    //: /sn:0 {0}(448,288)(448,208)(433,208)(433,177){1}
wire w9;    //: /sn:0 {0}(800,85)(800,296){1}
wire w51;    //: /sn:0 {0}(1066,511)(1066,622){1}
wire w57;    //: /sn:0 {0}(1036,511)(1036,622){1}
//: enddecls

  MUL4 g44 (.b(w45), .a(w46), .out(w47));   //: @(139, 388) /sz:(53, 56) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]
  assign w6 = b[1]; //: TAP g8 @(1051,171) /sn:0 /R:1 /w:[ 1 29 30 ] /ss:1
  assign w1 = a[1]; //: TAP g4 @(1093,79) /sn:0 /R:1 /w:[ 0 29 30 ] /ss:1
  assign w64 = {w40, w57, w53, w52, w51}; //: CONCAT g47  @(1046,627) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w9 = a[0]; //: TAP g16 @(800,79) /sn:0 /R:1 /w:[ 0 23 24 ] /ss:1
  assign w0 = a[0]; //: TAP g3 @(1107,79) /sn:0 /R:1 /w:[ 0 31 32 ] /ss:1
  assign w29 = a[6]; //: TAP g26 @(170,79) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w10 = a[1]; //: TAP g17 @(784,79) /sn:0 /R:1 /w:[ 0 21 22 ] /ss:1
  assign w2 = {w8, w7, w6, w5, w4, w3, w1, w0}; //: CONCAT g2  @(1072,293) /sn:0 /R:3 /w:[ 0 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  assign w26 = b[2]; //: TAP g30 @(433,171) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  assign w21 = a[4]; //: TAP g23 @(201,79) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  MUL4 g39 (.b(w37), .a(w36), .out(w54));   //: @(1045, 394) /sz:(53, 56) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]
  assign w22 = a[5]; //: TAP g24 @(185,79) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: IN g1 (b) @(1229,173) /sn:0 /R:2 /w:[ 33 ]
  //: GROUND g60 (w72) @(696,871) /sn:0 /R:1 /w:[ 0 ]
  assign w25 = b[0]; //: TAP g29 @(468,171) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  //: GROUND g51 (w40) @(1026,539) /sn:0 /R:2 /w:[ 0 ]
  assign w11 = a[2]; //: TAP g18 @(769,79) /sn:0 /R:1 /w:[ 1 19 20 ] /ss:1
  assign w28 = {w27, w26, w19, w25, w24, w23, w18, w20}; //: CONCAT g25  @(473,293) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  assign w8 = b[3]; //: TAP g10 @(1014,171) /sn:0 /R:1 /w:[ 1 25 26 ] /ss:1
  FA12 g64 (.b(w62), .a(w78), .cin(w72), .cout(w77), .s(w83));   //: @(578, 835) /sz:(77, 74) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  //: GROUND g49 (w58) @(709,700) /sn:0 /R:2 /w:[ 0 ]
  assign w68 = {w67, w66, w65, w63, w59}; //: CONCAT g50  @(447,637) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w4 = a[3]; //: TAP g6 @(1059,79) /sn:0 /R:1 /w:[ 1 25 26 ] /ss:1
  //: GROUND g58 (w71) @(218,705) /sn:0 /R:3 /w:[ 1 ]
  FA8 g56 (.a(w47), .b(w68), .cin(w70), .cout(w71), .s(w69));   //: @(261, 673) /sz:(69, 65) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w31 = a[7]; //: TAP g35 @(153,79) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w7 = b[2]; //: TAP g9 @(1032,171) /sn:0 /R:1 /w:[ 1 27 28 ] /ss:1
  assign w5 = b[0]; //: TAP g7 @(1067,171) /sn:0 /R:1 /w:[ 1 31 32 ] /ss:1
  assign w78 = {w69, w76, w75, w74, w73}; //: CONCAT g59  @(499,791) /sn:0 /R:3 /w:[ 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w30 = b[4]; //: TAP g31 @(161,171) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w20 = a[4]; //: TAP g22 @(508,79) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  //: GROUND g54 (w67) @(427,549) /sn:0 /R:2 /w:[ 0 ]
  assign {w42, w43} = w28; //: CONCAT g45  @(473,331) /sn:0 /R:1 /w:[ 0 0 0 ] /dr:0 /tp:0 /drp:0
  MUL4 g41 (.b(w38), .a(w39), .out(w41));   //: @(738, 395) /sz:(53, 56) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 ]
  assign w34 = b[7]; //: TAP g36 @(107,171) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w35 = {w34, w33, w32, w30, w31, w29, w22, w21}; //: CONCAT g33  @(166,301) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  FA8 g52 (.a(w41), .b(w64), .cin(w56), .cout(w60), .s(w61));   //: @(858, 662) /sz:(69, 65) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  assign {w45, w46} = w35; //: CONCAT g42  @(166,332) /sn:0 /R:1 /w:[ 0 0 0 ] /dr:0 /tp:0 /drp:0
  assign {w38, w39} = w17; //: CONCAT g40  @(765,339) /sn:0 /R:1 /w:[ 0 0 0 ] /dr:0 /tp:0 /drp:0
  assign w13 = b[4]; //: TAP g12 @(760,171) /sn:0 /R:1 /w:[ 1 23 24 ] /ss:1
  //: GROUND g57 (w70) @(365,704) /sn:0 /R:1 /w:[ 0 ]
  assign {w57, w53, w52, w51, w50, w55, w49, w48} = w54; //: CONCAT g46  @(1071,506) /sn:0 /R:1 /w:[ 0 0 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  assign w33 = b[6]; //: TAP g34 @(125,171) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w24 = a[7]; //: TAP g28 @(460,79) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign w15 = b[6]; //: TAP g14 @(724,171) /sn:0 /R:1 /w:[ 1 19 20 ] /ss:1
  assign w17 = {w16, w15, w14, w13, w12, w11, w10, w9}; //: CONCAT g11  @(765,301) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  assign w3 = a[2]; //: TAP g5 @(1077,79) /sn:0 /R:1 /w:[ 1 27 28 ] /ss:1
  //: GROUND g61 (w77) @(535,869) /sn:0 /R:3 /w:[ 0 ]
  assign w19 = b[1]; //: TAP g21 @(452,171) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  assign w12 = a[3]; //: TAP g19 @(752,79) /sn:0 /R:1 /w:[ 1 17 18 ] /ss:1
  assign w23 = a[6]; //: TAP g32 @(478,79) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  assign w18 = a[5]; //: TAP g20 @(494,79) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  //: OUT g63 (out) @(1095,1035) /sn:0 /R:3 /w:[ 1 ]
  MUL4 g43 (.b(w42), .a(w43), .out(w44));   //: @(446, 387) /sz:(53, 56) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]
  assign {w37, w36} = w2; //: CONCAT g38  @(1072,338) /sn:0 /R:1 /w:[ 0 0 1 ] /dr:0 /tp:0 /drp:0
  assign w16 = b[7]; //: TAP g15 @(706,171) /sn:0 /R:1 /w:[ 1 17 18 ] /ss:1
  //: IN g0 (a) @(1221,81) /sn:0 /R:2 /w:[ 33 ]
  assign w62 = {w58, w60, w61}; //: CONCAT g48  @(719,790) /sn:0 /R:3 /w:[ 1 1 1 0 ] /dr:1 /tp:0 /drp:1
  assign w27 = b[3]; //: TAP g27 @(415,171) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign out = {w83, w50, w55, w49, w48}; //: CONCAT g62  @(1095,995) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w32 = b[5]; //: TAP g37 @(145,171) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign {w66, w65, w63, w59, w76, w75, w74, w73} = w44; //: CONCAT g55  @(472,516) /sn:0 /R:1 /w:[ 0 0 0 0 0 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: GROUND g53 (w56) @(962,693) /sn:0 /R:1 /w:[ 0 ]
  assign w14 = b[5]; //: TAP g13 @(744,171) /sn:0 /R:1 /w:[ 1 21 22 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin MUL4
module MUL4(b, a, out);
//: interface  /sz:(56, 53) /bd:[ Li0>a[3:0](13/53) Li1>b[3:0](37/53) Ro0<out[7:0](26/53) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:638,-312)(567,-312){1}
//: {2}(566,-312)(426,-312){3}
//: {4}(425,-312)(368,-312){5}
//: {6}(367,-312)(54,-312){7}
//: {8}(53,-312)(46,-312){9}
supply0 w23;    //: /sn:0 {0}(88,79)(72,79){1}
supply0 w21;    //: /sn:0 {0}(311,91)(330,91){1}
output [7:0] out;    //: /sn:0 {0}(#:-133,771)(#:-133,809){1}
input [3:0] a;    //: /sn:0 {0}(#:-187,-180)(-180,-180){1}
//: {2}(-179,-180)(135,-180){3}
//: {4}(136,-180)(517,-180){5}
//: {6}(518,-180)(586,-180){7}
//: {8}(587,-180)(#:641,-180){9}
supply0 w9;    //: /sn:0 {0}(509,456)(516,456){1}
supply0 w26;    //: /sn:0 {0}(-139,537)(-123,537){1}
wire w16;    //: /sn:0 {0}(-578,252)(-578,215)(-520,215){1}
//: {2}(-516,215)(-409,215){3}
//: {4}(-407,213)(-407,-136)(-181,-136){5}
//: {6}(-179,-138)(-179,-176){7}
//: {8}(-179,-134)(-179,68){9}
//: {10}(-407,217)(-407,253){11}
//: {12}(-518,217)(-518,251){13}
wire w6;    //: /sn:0 {0}(498,-39)(498,-190)(565,-190){1}
//: {2}(567,-192)(567,-197){3}
//: {4}(567,-201)(567,-207){5}
//: {6}(567,-211)(567,-308){7}
//: {8}(565,-209)(-199,-209)(-199,68){9}
//: {10}(565,-199)(116,-199)(116,-44){11}
//: {12}(567,-188)(567,-39){13}
wire w13;    //: /sn:0 {0}(-148,765)(-148,676)(-384,676)(-384,566){1}
wire w7;    //: /sn:0 {0}(196,-44)(196,-87){1}
//: {2}(198,-89)(516,-89){3}
//: {4}(518,-91)(518,-100){5}
//: {6}(518,-104)(518,-176){7}
//: {8}(516,-102)(-245,-102)(-245,66){9}
//: {10}(518,-87)(518,-39){11}
//: {12}(194,-89)(-7,-89)(-7,-48){13}
wire w58;    //: /sn:0 {0}(-188,110)(-188,405)(-16,405)(-16,420){1}
wire w34;    //: /sn:0 {0}(136,-44)(136,-111){1}
//: {2}(136,-115)(136,-121){3}
//: {4}(136,-125)(136,-176){5}
//: {6}(134,-123)(-463,-123)(-463,254){7}
//: {8}(134,-113)(-113,-113)(-113,40){9}
//: {10}(-115,42)(-306,42)(-306,65){11}
//: {12}(-113,44)(-113,65){13}
wire w59;    //: /sn:0 {0}(-122,107)(-122,294)(3,294)(3,309){1}
wire w39;    //: /sn:0 {0}(34,454)(223,454){1}
wire w22;    //: /sn:0 {0}(509,3)(509,407)(490,407)(490,422){1}
wire w3;    //: /sn:0 {0}(426,-40)(426,-217){1}
//: {2}(426,-221)(426,-228){3}
//: {4}(426,-232)(426,-237){5}
//: {6}(426,-241)(426,-308){7}
//: {8}(424,-239)(-427,-239)(-427,253){9}
//: {10}(424,-230)(-133,-230)(-133,65){11}
//: {12}(424,-219)(176,-219)(176,-44){13}
wire w0;    //: /sn:0 {0}(368,-308)(368,-273){1}
//: {2}(366,-271)(-538,-271)(-538,251){3}
//: {4}(368,-269)(368,-261){5}
//: {6}(366,-259)(-326,-259)(-326,65){7}
//: {8}(368,-257)(368,-252){9}
//: {10}(366,-250)(13,-250)(13,-48){11}
//: {12}(368,-248)(368,-40){13}
wire w36;    //: /sn:0 {0}(-527,293)(-527,360)(-513,360)(-513,375){1}
wire w20;    //: /sn:0 {0}(65,-3)(65,30)(53,30)(53,45){1}
wire w60;    //: /sn:0 {0}(4,-6)(4,30)(22,30)(22,45){1}
wire w30;    //: /sn:0 {0}(-249,188)(-58,188)(-58,78)(3,78){1}
wire w29;    //: /sn:0 {0}(-35,453)(-158,453)(-158,503){1}
wire w37;    //: /sn:0 {0}(-287,218)(-287,308){1}
wire w42;    //: /sn:0 {0}(15,373)(15,420){1}
wire w18;    //: /sn:0 {0}(54,-45)(54,-277){1}
//: {2}(54,-281)(54,-286){3}
//: {4}(54,-290)(54,-308){5}
//: {6}(52,-288)(-483,-288)(-483,199){7}
//: {8}(-485,201)(-598,201)(-598,252){9}
//: {10}(-483,203)(-483,254){11}
//: {12}(52,-279)(-265,-279)(-265,66){13}
wire w12;    //: /sn:0 {0}(-138,765)(-138,663)(-177,663)(-177,567){1}
wire w19;    //: /sn:0 {0}(-168,765)(-168,701)(-621,701)(-621,534)(-606,534){1}
wire w10;    //: /sn:0 {0}(254,485)(254,668)(-118,668)(-118,765){1}
wire w54;    //: /sn:0 {0}(-537,535)(-415,535){1}
wire w24;    //: /sn:0 {0}(440,455)(292,455){1}
wire w1;    //: /sn:0 {0}(348,-40)(348,-66)(444,-66){1}
//: {2}(448,-66)(585,-66){3}
//: {4}(587,-68)(587,-74){5}
//: {6}(587,-78)(587,-176){7}
//: {8}(585,-76)(74,-76)(74,-45){9}
//: {10}(587,-64)(587,-39){11}
//: {12}(446,-64)(446,-40){13}
wire w31;    //: /sn:0 {0}(34,109)(34,309){1}
wire w8;    //: /sn:0 {0}(437,2)(437,407)(459,407)(459,422){1}
wire w46;    //: /sn:0 {0}(-416,295)(-416,298)(-318,298)(-318,308){1}
wire w17;    //: /sn:0 {0}(127,-2)(127,406)(242,406)(242,421){1}
wire w27;    //: /sn:0 {0}(242,90)(222,90)(222,343)(53,343){1}
wire w44;    //: /sn:0 {0}(-306,372)(-306,448)(-189,448)(-189,503){1}
wire w33;    //: /sn:0 {0}(-587,294)(-587,501){1}
wire w67;    //: /sn:0 {0}(-98,765)(-98,689)(578,689)(578,3){1}
wire w28;    //: /sn:0 {0}(273,121)(273,421){1}
wire w35;    //: /sn:0 {0}(-463,409)(-376,409)(-376,187)(-318,187){1}
wire w14;    //: /sn:0 {0}(187,-2)(187,42)(261,42)(261,57){1}
wire w45;    //: /sn:0 {0}(-532,408)(-556,408)(-556,501){1}
wire w2;    //: /sn:0 {0}(359,2)(359,42)(292,42)(292,57){1}
wire w48;    //: /sn:0 {0}(-315,107)(-315,139)(-299,139)(-299,154){1}
wire w11;    //: /sn:0 {0}(-128,765)(-128,654)(-4,654)(-4,484){1}
wire w41;    //: /sn:0 {0}(-16,342)(-268,342){1}
wire w47;    //: /sn:0 {0}(-501,439)(-501,487)(-396,487)(-396,502){1}
wire w15;    //: /sn:0 {0}(-158,765)(-158,688)(-575,688)(-575,565){1}
wire w38;    //: /sn:0 {0}(-472,296)(-472,360)(-482,360)(-482,375){1}
wire w5;    //: /sn:0 {0}(-108,765)(-108,680)(471,680)(471,486){1}
wire w43;    //: /sn:0 {0}(-337,341)(-365,341)(-365,502){1}
wire w57;    //: /sn:0 {0}(-254,108)(-254,139)(-268,139)(-268,154){1}
wire w51;    //: /sn:0 {0}(-346,536)(-208,536){1}
//: enddecls

  AND2 g4 (.in2(w6), .in1(w1), .out(w67));   //: @(557, -38) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>11 Bo0<1 ]
  AND2 g8 (.in2(w7), .in1(w0), .out(w60));   //: @(-17, -47) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>11 Bo0<0 ]
  //: joint g44 (w0) @(368, -259) /w:[ -1 5 6 8 ]
  AND2 g3 (.in2(w6), .in1(w7), .out(w22));   //: @(488, -38) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>11 Bo0<0 ]
  AND2 g16 (.in2(w3), .in1(w16), .out(w46));   //: @(-437, 254) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>9 Ti1>11 Bo0<0 ]
  //: joint g47 (w18) @(54, -279) /w:[ -1 2 12 1 ]
  //: IN g17 (b) @(640,-312) /sn:0 /R:2 /w:[ 0 ]
  assign w34 = a[2]; //: TAP g26 @(136,-182) /sn:0 /R:1 /w:[ 5 3 4 ] /ss:1
  AND2 g2 (.in2(w3), .in1(w1), .out(w8));   //: @(416, -39) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>13 Bo0<0 ]
  //: joint g23 (w7) @(518, -89) /w:[ -1 4 3 10 ]
  assign w16 = a[3]; //: TAP g30 @(-179,-182) /sn:0 /R:1 /w:[ 7 1 2 ] /ss:1
  //: IN g1 (a) @(643,-180) /sn:0 /R:2 /w:[ 9 ]
  //: joint g24 (w7) @(196, -89) /w:[ 2 -1 12 1 ]
  //: joint g39 (w3) @(426, -219) /w:[ -1 2 12 1 ]
  //: joint g29 (w34) @(136, -123) /w:[ -1 4 6 3 ]
  FA2 g60 (.b(w37), .a(w46), .cin(w41), .cout(w43), .s(w44));   //: @(-336, 309) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA2 g51 (.b(w22), .a(w8), .cin(w9), .cout(w24), .s(w5));   //: @(441, 423) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<1 ]
  assign w1 = a[0]; //: TAP g18 @(587,-182) /sn:0 /R:1 /w:[ 7 7 8 ] /ss:1
  AND2 g10 (.in2(w6), .in1(w16), .out(w58));   //: @(-209, 69) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>9 Ti1>9 Bo0<0 ]
  //: joint g25 (w7) @(518, -102) /w:[ -1 6 8 5 ]
  FA2 g65 (.b(w43), .a(w47), .cin(w51), .cout(w54), .s(w13));   //: @(-414, 503) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  //: GROUND g64 (w26) @(-117,537) /sn:0 /R:1 /w:[ 1 ]
  //: joint g49 (w18) @(-483, 201) /w:[ -1 7 8 10 ]
  AND2 g6 (.in2(w6), .in1(w34), .out(w17));   //: @(106, -43) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>11 Ti1>0 Bo0<0 ]
  assign out = {w19, w15, w13, w12, w11, w10, w5, w67}; //: CONCAT g50  @(-133,770) /sn:0 /R:3 /w:[ 0 0 0 0 0 0 1 0 0 ] /dr:1 /tp:0 /drp:1
  //: OUT g68 (out) @(-133,806) /sn:0 /R:3 /w:[ 1 ]
  AND2 g7 (.in2(w18), .in1(w1), .out(w20));   //: @(44, -44) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>9 Bo0<0 ]
  AND2 g9 (.in2(w3), .in1(w34), .out(w59));   //: @(-143, 66) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>11 Ti1>13 Bo0<0 ]
  //: joint g35 (w6) @(567, -190) /w:[ -1 2 1 12 ]
  FA2 g56 (.b(w57), .a(w48), .cin(w30), .cout(w35), .s(w37));   //: @(-317, 155) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  FA2 g58 (.b(w28), .a(w17), .cin(w24), .cout(w39), .s(w10));   //: @(224, 422) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  //: joint g22 (w1) @(587, -76) /w:[ -1 6 8 5 ]
  //: joint g31 (w16) @(-179, -136) /w:[ -1 6 5 8 ]
  FA2 g59 (.b(w31), .a(w59), .cin(w27), .cout(w41), .s(w42));   //: @(-15, 310) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g33 (w16) @(-407, 215) /w:[ -1 4 3 10 ]
  //: joint g36 (w6) @(567, -199) /w:[ -1 4 10 3 ]
  //: joint g41 (w3) @(426, -239) /w:[ -1 6 8 5 ]
  //: joint g45 (w0) @(368, -271) /w:[ -1 1 2 4 ]
  //: GROUND g54 (w21) @(336,91) /sn:0 /R:1 /w:[ 1 ]
  //: joint g40 (w3) @(426, -230) /w:[ -1 4 10 3 ]
  assign w0 = b[2]; //: TAP g42 @(368,-314) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: GROUND g52 (w9) @(522,456) /sn:0 /R:1 /w:[ 1 ]
  FA2 g66 (.b(w45), .a(w33), .cin(w54), .cout(w19), .s(w15));   //: @(-605, 502) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  AND2 g12 (.in2(w0), .in1(w34), .out(w48));   //: @(-336, 66) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>7 Ti1>11 Bo0<0 ]
  //: joint g28 (w34) @(-113, 42) /w:[ -1 9 10 12 ]
  assign w6 = b[0]; //: TAP g34 @(567,-314) /sn:0 /R:1 /w:[ 7 2 1 ] /ss:1
  assign w18 = b[3]; //: TAP g46 @(54,-314) /sn:0 /R:1 /w:[ 5 8 7 ] /ss:1
  //: GROUND g57 (w23) @(94,79) /sn:0 /R:1 /w:[ 0 ]
  AND2 g5 (.in2(w3), .in1(w7), .out(w14));   //: @(166, -43) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>0 Bo0<0 ]
  AND2 g11 (.in2(w18), .in1(w7), .out(w57));   //: @(-275, 67) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>13 Ti1>9 Bo0<0 ]
  AND2 g14 (.in2(w0), .in1(w16), .out(w36));   //: @(-548, 252) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>3 Ti1>13 Bo0<0 ]
  assign w7 = a[1]; //: TAP g21 @(518,-182) /sn:0 /R:1 /w:[ 7 5 6 ] /ss:1
  //: joint g19 (w1) @(587, -66) /w:[ -1 4 3 10 ]
  FA2 g61 (.b(w38), .a(w36), .cin(w35), .cout(w45), .s(w47));   //: @(-531, 376) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g32 (w16) @(-518, 215) /w:[ 2 -1 1 12 ]
  //: joint g20 (w1) @(446, -66) /w:[ 2 -1 1 12 ]
  FA2 g63 (.b(w29), .a(w44), .cin(w26), .cout(w51), .s(w12));   //: @(-207, 504) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  AND2 g0 (.in2(w1), .in1(w0), .out(w2));   //: @(338, -39) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>0 Ti1>13 Bo0<0 ]
  AND2 g15 (.in2(w18), .in1(w34), .out(w38));   //: @(-493, 255) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>11 Ti1>7 Bo0<0 ]
  assign w3 = b[1]; //: TAP g38 @(426,-314) /sn:0 /R:1 /w:[ 7 4 3 ] /ss:1
  //: joint g43 (w0) @(368, -250) /w:[ -1 9 10 12 ]
  //: joint g27 (w34) @(136, -113) /w:[ -1 2 8 1 ]
  //: joint g48 (w18) @(54, -288) /w:[ -1 4 6 3 ]
  //: joint g37 (w6) @(567, -209) /w:[ -1 6 8 5 ]
  FA2 g62 (.b(w42), .a(w58), .cin(w39), .cout(w29), .s(w11));   //: @(-34, 421) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<1 ]
  FA2 g55 (.b(w20), .a(w60), .cin(w23), .cout(w30), .s(w31));   //: @(4, 46) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  AND2 g13 (.in2(w18), .in1(w16), .out(w33));   //: @(-608, 253) /sz:(40, 40) /R:3 /sn:0 /p:[ Ti0>9 Ti1>0 Bo0<0 ]
  FA2 g53 (.b(w2), .a(w14), .cin(w21), .cout(w27), .s(w28));   //: @(243, 58) /sz:(67, 62) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA8
module FA8(b, cin, cout, a, s);
//: interface  /sz:(69, 65) /bd:[ Ti0>b[7:0](47/69) Ti1>a[7:0](14/69) Ri0>cin(31/65) Lo0<cout(32/65) Bo0<s[7:0](32/69) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [7:0] b;    //: /sn:0 {0}(#:250,167)(258,167){1}
//: {2}(259,167)(271,167){3}
//: {4}(272,167)(286,167){5}
//: {6}(287,167)(301,167){7}
//: {8}(302,167)(451,167){9}
//: {10}(452,167)(468,167){11}
//: {12}(469,167)(488,167){13}
//: {14}(489,167)(505,167){15}
//: {16}(506,167)(#:707,167){17}
input cin;    //: /sn:0 {0}(534,353)(573,353){1}
output cout;    //: /sn:0 {0}(288,353)(266,353)(266,485){1}
output [7:0] s;    //: /sn:0 {0}(402,492)(#:402,439){1}
input [7:0] a;    //: /sn:0 {0}(#:704,107)(568,107){1}
//: {2}(567,107)(551,107){3}
//: {4}(550,107)(535,107){5}
//: {6}(534,107)(516,107){7}
//: {8}(515,107)(355,107){9}
//: {10}(354,107)(340,107){11}
//: {12}(339,107)(325,107){13}
//: {14}(324,107)(312,107){15}
//: {16}(311,107)(303,107){17}
wire w6;    //: /sn:0 {0}(292,233)(292,196)(287,196)(287,171){1}
wire w13;    //: /sn:0 {0}(506,237)(506,171){1}
wire w16;    //: /sn:0 {0}(476,237)(476,219)(452,219)(452,171){1}
wire w7;    //: /sn:0 {0}(282,233)(282,204)(272,204)(272,171){1}
wire w4;    //: /sn:0 {0}(312,233)(312,111){1}
wire [3:0] w22;    //: /sn:0 {0}(#:299,333)(299,305)(302,305)(302,289){1}
wire w0;    //: /sn:0 {0}(355,111)(355,214)(342,214)(342,233){1}
wire w3;    //: /sn:0 {0}(322,233)(322,194)(325,194)(325,111){1}
wire [3:0] w20;    //: /sn:0 {0}(#:521,333)(521,310)(516,310)(516,288){1}
wire w18;    //: /sn:0 {0}(492,353)(330,353){1}
wire w12;    //: /sn:0 {0}(516,237)(516,111){1}
wire [3:0] w19;    //: /sn:0 {0}(#:397,433)(397,401)(306,401)(#:306,375){1}
wire [3:0] w23;    //: /sn:0 {0}(#:317,333)(317,306)(312,306)(312,289){1}
wire w10;    //: /sn:0 {0}(551,111)(551,204)(536,204)(536,237){1}
wire [3:0] w24;    //: /sn:0 {0}(407,433)(407,401)(#:510,401)(#:510,375){1}
wire [3:0] w21;    //: /sn:0 {0}(#:503,333)(503,308)(506,308)(506,288){1}
wire w1;    //: /sn:0 {0}(340,111)(340,203)(332,203)(332,233){1}
wire w8;    //: /sn:0 {0}(272,233)(272,212)(259,212)(259,171){1}
wire [7:0] w17;    //: /sn:0 {0}(#:511,282)(#:511,243){1}
wire w14;    //: /sn:0 {0}(496,237)(496,193)(489,193)(489,171){1}
wire [7:0] w2;    //: /sn:0 {0}(#:307,239)(#:307,283){1}
wire w11;    //: /sn:0 {0}(526,237)(526,190)(535,190)(535,111){1}
wire w15;    //: /sn:0 {0}(486,237)(486,206)(469,206)(469,171){1}
wire w5;    //: /sn:0 {0}(302,233)(302,171){1}
wire w9;    //: /sn:0 {0}(568,111)(568,216)(546,216)(546,237){1}
//: enddecls

  assign w9 = a[0]; //: TAP g4 @(568,105) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  assign w13 = b[0]; //: TAP g8 @(506,165) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  assign w17 = {w16, w15, w14, w13, w12, w11, w10, w9}; //: CONCAT g3  @(511,242) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  assign w5 = b[4]; //: TAP g16 @(302,165) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w6 = b[5]; //: TAP g17 @(287,165) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign s = {w19, w24}; //: CONCAT g26  @(402,438) /sn:0 /R:3 /w:[ 1 0 0 ] /dr:1 /tp:0 /drp:1
  assign w2 = {w8, w7, w6, w5, w4, w3, w1, w0}; //: CONCAT g2  @(307,238) /sn:0 /R:3 /w:[ 0 0 0 0 0 0 0 1 1 ] /dr:1 /tp:0 /drp:1
  FA4 g23 (.a(w21), .b(w20), .cin(cin), .cout(w18), .s(w24));   //: @(493, 334) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  //: IN g1 (b) @(709,167) /sn:0 /R:2 /w:[ 17 ]
  //: IN g24 (cin) @(575,353) /sn:0 /R:2 /w:[ 1 ]
  assign w7 = b[6]; //: TAP g18 @(272,165) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w15 = b[2]; //: TAP g10 @(469,165) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  //: OUT g25 (cout) @(266,482) /sn:0 /R:3 /w:[ 1 ]
  assign w11 = a[2]; //: TAP g6 @(535,105) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  assign w12 = a[3]; //: TAP g7 @(516,105) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  assign w14 = b[1]; //: TAP g9 @(489,165) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  FA4 g22 (.a(w22), .b(w23), .cin(w18), .cout(cout), .s(w19));   //: @(289, 334) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w0 = a[4]; //: TAP g12 @(355,105) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  assign w10 = a[1]; //: TAP g5 @(551,105) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  assign w16 = b[3]; //: TAP g11 @(452,165) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign w3 = a[6]; //: TAP g14 @(325,105) /sn:0 /R:1 /w:[ 1 14 13 ] /ss:1
  assign w8 = b[7]; //: TAP g19 @(259,165) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign {w21, w20} = w17; //: CONCAT g21  @(511,283) /sn:0 /R:1 /w:[ 1 1 0 ] /dr:0 /tp:0 /drp:0
  assign {w22, w23} = w2; //: CONCAT g20  @(307,284) /sn:0 /R:1 /w:[ 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: IN g0 (a) @(706,107) /sn:0 /R:2 /w:[ 0 ]
  assign w4 = a[7]; //: TAP g15 @(312,105) /sn:0 /R:1 /w:[ 1 16 15 ] /ss:1
  //: OUT g27 (s) @(402,489) /sn:0 /R:3 /w:[ 0 ]
  assign w1 = a[5]; //: TAP g13 @(340,105) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin REG16
module REG16(clk, out, in);
//: interface  /sz:(64, 59) /bd:[ Li0>in[15:0](29/59) Bi0>clk(32/64) Ro0<out[15:0](29/59) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [15:0] in;    //: /sn:0 {0}(#:725,539)(725,531){1}
//: {2}(725,530)(725,457){3}
//: {4}(725,456)(725,382){5}
//: {6}(725,381)(725,310){7}
//: {8}(725,309)(725,242){9}
//: {10}(725,241)(725,175){11}
//: {12}(725,174)(725,103){13}
//: {14}(725,102)(725,40){15}
//: {16}(725,39)(725,-5)(193,-5){17}
//: {18}(189,-5)(#:142,-5){19}
//: {20}(191,-3)(191,35){21}
//: {22}(191,36)(191,109){23}
//: {24}(191,110)(191,184){25}
//: {26}(191,185)(191,256){27}
//: {28}(191,257)(191,324){29}
//: {30}(191,325)(191,391){31}
//: {32}(191,392)(191,463){33}
//: {34}(191,464)(191,526){35}
//: {36}(191,527)(191,534){37}
input clk;    //: /sn:0 {0}(613,508)(613,490)(670,490)(670,418){1}
//: {2}(668,416)(615,416)(615,434){3}
//: {4}(670,414)(670,341){5}
//: {6}(668,339)(614,339)(614,359){7}
//: {8}(670,337)(670,271){9}
//: {10}(668,269)(614,269)(614,287){11}
//: {12}(670,267)(670,215){13}
//: {14}(668,213)(614,213)(614,219){15}
//: {16}(670,211)(670,144){17}
//: {18}(668,142)(616,142)(616,152){19}
//: {20}(670,140)(670,69){21}
//: {22}(670,65)(670,7){23}
//: {24}(670,3)(670,-23)(247,-23)(247,74){25}
//: {26}(249,76)(304,76)(304,58){27}
//: {28}(247,78)(247,148){29}
//: {30}(249,150)(302,150)(302,132){31}
//: {32}(247,152)(247,225){33}
//: {34}(249,227)(303,227)(303,207){35}
//: {36}(247,229)(247,295){37}
//: {38}(249,297)(303,297)(303,279){39}
//: {40}(247,299)(247,351){41}
//: {42}(249,353)(303,353)(303,347){43}
//: {44}(245,353)(146,353){45}
//: {46}(247,355)(247,422){47}
//: {48}(249,424)(301,424)(301,414){49}
//: {50}(247,426)(247,497){51}
//: {52}(249,499)(298,499)(298,486){53}
//: {54}(247,501)(247,561)(297,561)(297,549){55}
//: {56}(668,5)(620,5)(620,17){57}
//: {58}(668,67)(619,67)(619,80){59}
output [15:0] out;    //: /sn:0 {0}(#:463,630)(463,688)(462,688)(462,692){1}
wire w6;    //: /sn:0 {0}(195,185)(284,185){1}
wire w13;    //: /sn:0 {0}(591,309)(508,309)(508,624){1}
wire w16;    //: /sn:0 {0}(591,381)(518,381)(518,624){1}
wire w7;    //: /sn:0 {0}(593,174)(488,174)(488,624){1}
wire w4;    //: /sn:0 {0}(325,110)(398,110)(398,624){1}
wire w3;    //: /sn:0 {0}(195,110)(283,110){1}
wire w0;    //: /sn:0 {0}(195,36)(285,36){1}
wire w22;    //: /sn:0 {0}(590,530)(538,530)(538,624){1}
wire w36;    //: /sn:0 {0}(730,174)(635,174){1}
wire w20;    //: /sn:0 {0}(321,464)(448,464)(448,624){1}
wire w30;    //: /sn:0 {0}(730,102)(638,102){1}
wire w18;    //: /sn:0 {0}(195,464)(279,464){1}
wire w12;    //: /sn:0 {0}(195,392)(282,392){1}
wire w19;    //: /sn:0 {0}(592,456)(528,456)(528,624){1}
wire w23;    //: /sn:0 {0}(320,527)(458,527)(458,624){1}
wire w10;    //: /sn:0 {0}(591,241)(498,241)(498,624){1}
wire w21;    //: /sn:0 {0}(195,527)(278,527){1}
wire w24;    //: /sn:0 {0}(730,241)(633,241){1}
wire w1;    //: /sn:0 {0}(468,624)(468,39)(597,39){1}
wire w31;    //: /sn:0 {0}(730,39)(639,39){1}
wire w8;    //: /sn:0 {0}(326,185)(408,185)(408,624){1}
wire w17;    //: /sn:0 {0}(326,325)(428,325)(428,624){1}
wire w28;    //: /sn:0 {0}(730,530)(632,530){1}
wire w33;    //: /sn:0 {0}(730,309)(633,309){1}
wire w14;    //: /sn:0 {0}(324,392)(438,392)(438,624){1}
wire w11;    //: /sn:0 {0}(326,257)(418,257)(418,624){1}
wire w2;    //: /sn:0 {0}(327,36)(388,36)(388,624){1}
wire w15;    //: /sn:0 {0}(195,325)(284,325){1}
wire w5;    //: /sn:0 {0}(596,102)(478,102)(478,624){1}
wire w38;    //: /sn:0 {0}(730,381)(633,381){1}
wire w9;    //: /sn:0 {0}(195,257)(284,257){1}
wire w26;    //: /sn:0 {0}(730,456)(634,456){1}
//: enddecls

  FFD g8 (.D(w15), .Clk(clk), .Y(w17));   //: @(285, 306) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>43 Ro0<0 ]
  FFD g4 (.D(w3), .Clk(clk), .Y(w4));   //: @(284, 91) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>31 Ro0<0 ]
  FFD g44 (.Clk(clk), .D(w38), .Y(w16));   //: @(592, 360) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>7 Ri0>1 Lo0<0 ]
  FFD g3 (.D(w0), .Clk(clk), .Y(w2));   //: @(286, 17) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>27 Ro0<0 ]
  //: joint g16 (clk) @(247, 499) /w:[ 52 51 -1 54 ]
  //: joint g47 (clk) @(670, 142) /w:[ 18 17 -1 20 ]
  assign w0 = in[0]; //: TAP g17 @(189,36) /sn:0 /R:2 /w:[ 0 22 21 ] /ss:1
  //: joint g26 (clk) @(670, 67) /w:[ -1 22 58 21 ]
  //: IN g2 (clk) @(144,353) /sn:0 /w:[ 45 ]
  assign w18 = in[6]; //: TAP g23 @(189,464) /sn:0 /R:2 /w:[ 0 34 33 ] /ss:1
  assign w28 = in[15]; //: TAP g30 @(728,530) /sn:0 /w:[ 0 2 1 ] /ss:1
  //: OUT g1 (out) @(462,689) /sn:0 /R:3 /w:[ 1 ]
  assign w21 = in[7]; //: TAP g24 @(189,527) /sn:0 /R:2 /w:[ 0 36 35 ] /ss:1
  FFD g39 (.Clk(clk), .D(w36), .Y(w7));   //: @(594, 153) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>19 Ri0>1 Lo0<0 ]
  FFD g29 (.Clk(clk), .D(w28), .Y(w22));   //: @(591, 509) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>0 Ri0>1 Lo0<0 ]
  assign w3 = in[1]; //: TAP g18 @(189,110) /sn:0 /R:2 /w:[ 0 24 23 ] /ss:1
  FFD g10 (.D(w21), .Clk(clk), .Y(w23));   //: @(279, 508) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>55 Ro0<0 ]
  assign out = {w22, w19, w16, w13, w10, w7, w5, w1, w23, w20, w14, w17, w11, w8, w4, w2}; //: CONCAT g25  @(463,629) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  //: joint g49 (clk) @(670, 269) /w:[ 10 9 -1 12 ]
  FFD g6 (.D(w9), .Clk(clk), .Y(w11));   //: @(285, 238) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>39 Ro0<0 ]
  //: joint g50 (clk) @(670, 5) /w:[ -1 24 56 23 ]
  FFD g9 (.D(w18), .Clk(clk), .Y(w20));   //: @(280, 445) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>53 Ro0<0 ]
  FFD g7 (.D(w12), .Clk(clk), .Y(w14));   //: @(283, 373) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>49 Ro0<0 ]
  assign w36 = in[10]; //: TAP g35 @(728,174) /sn:0 /w:[ 0 12 11 ] /ss:1
  assign w12 = in[5]; //: TAP g22 @(189,392) /sn:0 /R:2 /w:[ 0 32 31 ] /ss:1
  //: joint g31 (clk) @(247, 76) /w:[ 26 25 -1 28 ]
  assign w31 = in[8]; //: TAP g33 @(728,39) /sn:0 /w:[ 0 16 15 ] /ss:1
  FFD g36 (.Clk(clk), .D(w31), .Y(w1));   //: @(598, 18) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>57 Ri0>1 Lo0<1 ]
  //: joint g41 (clk) @(670, 416) /w:[ 2 1 -1 4 ]
  assign w24 = in[11]; //: TAP g45 @(728,241) /sn:0 /w:[ 0 10 9 ] /ss:1
  //: joint g40 (clk) @(670, 339) /w:[ 6 5 -1 8 ]
  //: joint g42 (clk) @(670, 213) /w:[ 14 13 -1 16 ]
  //: joint g12 (clk) @(247, 227) /w:[ 34 33 -1 36 ]
  FFD g28 (.Clk(clk), .D(w26), .Y(w19));   //: @(593, 435) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>3 Ri0>1 Lo0<0 ]
  assign w26 = in[14]; //: TAP g34 @(728,456) /sn:0 /w:[ 0 4 3 ] /ss:1
  assign w33 = in[12]; //: TAP g46 @(728,309) /sn:0 /w:[ 0 8 7 ] /ss:1
  //: joint g11 (clk) @(247, 150) /w:[ 30 29 -1 32 ]
  //: joint g14 (clk) @(247, 353) /w:[ 42 41 44 46 ]
  FFD g5 (.D(w6), .Clk(clk), .Y(w8));   //: @(285, 166) /sz:(40, 40) /sn:0 /p:[ Li0>1 Bi0>35 Ro0<0 ]
  assign w6 = in[2]; //: TAP g19 @(189,185) /sn:0 /R:2 /w:[ 0 26 25 ] /ss:1
  assign w15 = in[4]; //: TAP g21 @(189,325) /sn:0 /R:2 /w:[ 0 30 29 ] /ss:1
  assign w9 = in[3]; //: TAP g20 @(189,257) /sn:0 /R:2 /w:[ 0 28 27 ] /ss:1
  assign w30 = in[9]; //: TAP g32 @(728,102) /sn:0 /w:[ 0 14 13 ] /ss:1
  //: joint g15 (clk) @(247, 424) /w:[ 48 47 -1 50 ]
  //: IN g0 (in) @(140,-5) /sn:0 /w:[ 19 ]
  FFD g38 (.Clk(clk), .D(w30), .Y(w5));   //: @(597, 81) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>59 Ri0>1 Lo0<0 ]
  assign w38 = in[13]; //: TAP g43 @(728,381) /sn:0 /w:[ 0 6 5 ] /ss:1
  FFD g27 (.Clk(clk), .D(w24), .Y(w10));   //: @(592, 220) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>15 Ri0>1 Lo0<0 ]
  //: joint g48 (in) @(191, -5) /w:[ 17 -1 18 20 ]
  FFD g37 (.Clk(clk), .D(w33), .Y(w13));   //: @(592, 288) /sz:(40, 40) /R:2 /sn:0 /p:[ Ti0>11 Ri0>1 Lo0<0 ]
  //: joint g13 (clk) @(247, 297) /w:[ 38 37 -1 40 ]

endmodule
//: /netlistEnd

